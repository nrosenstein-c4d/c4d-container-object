MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ����mǉ�mǉ�mǉ~��mǉ�mƉ�mǉ���mǉd� ��mǉ�
��mǉ�	��mǉ���mǉa���mǉa���mǉa���mǉRich�mǉ        PE  d� i{�Q        � "     D     ��       �                        �         `                                   �� ^   ` <            � �\           p �   ( 8                           @S p           �b �                          .text   j                        `.rdata  >�      �   
             @  @.data   q   �     �             @  �.pdata  g   �  h   �             @  @.idata  �	   `  
   4             @  �.reloc  �   p     >             @  B                                                                                                                                                                                                                                                                                        ������6  ��	  ��  �W  �R  ��  ��  ��  ��  �I  �  �o  ��  �  �0  �	  �  �A  ��  ��  �B	  ��  �H  �
  �
  �9  �  ��  ��  ��  ��  ��  �  �	  ��  �  ��  �-  ��  �  �^  �I  �  �  �J  ��  �   �k  �  �  �  ��  ��  �=	  ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������H��(�I����   H��(������������������������������H�T$�L$H��8�D$@�D$ �|$ t�H��� ��   ��   H��8���������������������������H�L$H��(A�E3�3�H�L$0��  H��(�����������������H�L$H��(H�L$0�}  H��(���������L�L$ D�D$H�T$H�L$H��(�D$@�ȉD$@�|$@ | H�L$0�T$HH�D$8H�L$0H�H��H�D$0��H��(�����������������������������������D�L$ D�D$�T$H�L$H��H�D$0    �H�L$P����H�D$PH�|$P t{D�D$`�T$XH�L$P�5y  H�L$P�Y���H�D$8�|$h tCH�|$8 t;�D$     D�L$hD�D$`�T$XH�L$8�����D$4�|$p t�D$4�L$0ȋ��D$0�D$0���D$0�n����D$0H��H���������������������D�L$ D�D$�T$H�L$H��8�D$     �H�L$@�����H�D$@H�|$@ t1�T$HH�L$@�*x  �D$$�D$P9D$$u�D$ ���D$ �|$X t�븋D$ H��8���������������H��   H�D$`����E3�H�� H�L$h������H�T$hH�L$H�L�  �H�L$h������D$X    �D$\    E3�H�� H��$�   �����H�L$H�`���H�D$P3��!  �D$0    H�L$PH�L$(H��$�   H�L$ L����E3�H�йD� �� �D$@H��$�   �g����H�L$H衊  �D$@H�Ĩ   ������������������������������������������������������������������������������������������������������������������������������������������������������H�L$H��(H�L$0����H�D$0H�� H�H�D$0H��(����������������������\$ �T$�L$H�L$H�D$�D$� H�D$�D$�@H�D$�D$ �@H�D$���������������������H�L$H�D$W�� H�D$W��@H�D$W��@H�D$����������������H�L$H��(H�L$0�2  H�D$0H�� H�H�D$0H��(���������������������H�L$H��(H�L$0�����H�D$0H�) H�H�D$0H��(���������������������H�T$H�L$H��(H��� H�@(H�L$0�PH��� H�@(H�T$0H�L$8�P8H�D$0H��(������������������������������D�D$H�T$H�L$H��(H�n� H�@(H�L$0�PH�[� H�@(D�L$@A�����H�T$8H�L$0�P H�D$0H��(������������������������������H�L$H��(H�� H�@(H�L$0�PH�D$0H��(�����������H�L$H��(H�L$0�a���H��(���������H�L$H��(H�L$0�0  H��(���������H�L$H��(H�L$0�����H��(���������H�L$H��(H�x� H�@(H�L$0�P0H��(����������������L�L$ D�D$H�T$H�L$H��(A�L�D$H�T$@H�L$0�R  H��(��������������L�L$ D�D$H�T$H�L$H��(H�L$0��  H��(����������H�L$H�D$H� ������������������̉T$H�L$H��(H�L$0�8����D$8����t
H�L$0�
���H�D$0H��(��������������������������̉T$H�L$H��(H�L$0�����D$8����t
H�L$0����H�D$0H��(��������������������������̉T$H�L$H��(H�L$0�����D$8����t
H�L$0�j���H�D$0H��(���������������������������H��HH�D$8����L�t A�E   H��� �   ����H�D$ H�|$  tH�L$ �����H�D$(�	H�D$(    H�D$(H�D$0H�D$0H��H���������������������������L�L$ L�D$H�T$H�L$H��HH�D$xH�D$(�D$p�D$ L�L$hL�D$`H�T$XH�L$P�  �D$0�|$0 u�D$0�BH�D$XH�D$8H�D$8H�x tH�D$8H��H��赒  H�D$PH�H��  H�L$8H�A�D$0H��H������������������������������������������������������H�T$H�L$H��(H�T$8H�L$0��}  H�D$0H�x tH�D$0H��H���&�  H��(������������������H�L$H��(H�(� H�@0H�L$0�P H��(����������������H�L$H��(H��� H�@0H�L$0�PH��(����������������H�L$H��(H��� H���   H�L$0�PXH��(�������������H�L$H��(H��� H��  H�L$0�PhH��(�������������H�L$H��(H�h� H��  H�L$0�PhH��(�������������D�D$�T$H�L$H��(H�/� H�@ D�D$@�T$8H�L$0��@  H��(���������������������������H�L$H��(H��� H��  H�L$0�PPH��(�������������L�L$ D�D$H�T$H�L$VWH��HH��� H�@ L�L$xD�D$pH�T$ H�L$`��`  H�|$hH��   �H�D$hH��H_^�����������������������H�T$H�L$H��XH�T$hH�L$`�{  �D$ �|$  u�D$ �yH�L$h�k���H�D$(A�   ��  H�L$(������� �� �� H�L$0� ���L����  H�L$(�s���H�D$`H�x tH�D$`H��H��荏  �D$ H��X����������������������������������������������������̉T$H�L$H��hH�D$8�����D$     H�S� H�@(�T$xH�L$@�PPH�D$(H�D$(H�D$0H�T$0H�L$p�M����D$ ���D$ H�L$@����H�D$pH��h�������������������������������L�L$ D�D$H�T$H�L$H��8L�L$XD�D$PH�T$HH�L$@�z  �D$$�|$$ u�D$$�kH�D$HH�D$(�D$P�D$ �|$ t�|$ t"�|$ �F t)�;L�D$XH�T$(H�L$@�����%H�T$(H�L$@�d����L�D$XH�T$(H�L$@�!����D$$H��8�����������������������������������������������L�D$H�T$H�L$H��  HǄ$�   ����H��$0  H���^� ��H��$0  ���� � �D$<�D$0�����D$<�D$4�D$4-�  �D$4�|$4�)  HcD$4H�������l$  H���H��$(  �V �D$     A�   A�   �?   H��������D$8�D$0�  ��  �D$8    H��$(  �SV �D$     A�   A�   �?   H�������D$0�  �  H��$(  �����D$     A�   A�   �?   H���k����D$8�D$0�  �P  �D$8    H��$(  �:����D$     A�   A�   �?   H���$����D$0�  �  H��$�   �+  ��   H��$�   ��c  H��$�   H��$�   H�D$`H�T$`H��$�   �L1  �H��$�   ��,  H��$�   ����H�D$PH�D$PH�D$x�   �H  H�L$xH�L$ L��E3��   H��$�   �6-  �D$DH��$�   �@����|$D �"  H��$   H�x u�f�  H��$   H�A�H��$   H�H臄  H��$   H�x u�   �  H���&% ��   E3�A�����H��$�   H��$   H�H�?�  �D$@�|$@t �   �% H��$   H��H�����  �|�ϊ  H�D$H�D$     A�   A�@   �@   H�L$H�7�  �D$    A�   A�   H�T$HH��$   H�H���  H��$   H��H��艊  H��$   H�L$HH�HH��$�   �[+  �#H��$   H�x tH��$   H��H���F�  �|$0 |SH��$(  ����H�D$X�T$8H��$�   �����H�D$hH�D$hH�D$pL�D$p�T$0H�L$X�w����H��$�   ����H��  �{!  �!  
$  �   8!  
$  
$  �!  �#  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L�D$H�T$H�L$H���   H��$�   H� H�D$8H��$�   H�x twH�D$8H�8 t%H�D$8H� H�D$0H�T$0H��$�   H�H�-�  �H��$�   H�H蚀  H�D$0�D$d    �D$h    H�L$0�W����D$HH�L$0�!����D$T�   H�D$8H� H�D$0H�|$0 u-�ʇ  H�D$0�D$     A�   A�@   �@   H�L$0�2�  H�T$8�D� �� ��tH�T$0H�D$8H��}�  H�D$8�@�D$dH�D$8�@�D$hH�D$8�@�D$HH�D$8�@�D$TH�|$0 ��  H��$�   �����H��$�   E3���  H��$�   �����D$L�|$L �i  H��$�   ����L��A��  H��$�   H��$�   ������ �Y�$�   �,��D$p� �Y�$�   �,��D$t�� �Y�$�   �,��D$lH�L$0藄  H�D$x�D$H�������D$L�D$LH��$�   �8���A�   A�   �?   H����������   �D$X    �
�D$X���D$X�D$H9D$X��   �D$X�D$@�D$P   �
�D$P���D$P�D$L9D$Pg�D$T�L$hȋ�+D$P�D$D�D$l�D$(�D$t�D$ D�L$pD�D$D�T$@H�L$0�����H�|$x t!�D$ �   D�L$DD�D$@H�T$xH�L$0������V���H��$�   ��N A�   A�   �?   H���9�������   �D$`    �
�D$`���D$`�D$T9D$`��   �D$`�D$D�D$\   �
�D$\���D$\�D$L9D$\g�D$H�L$dȋ�+D$\�D$@�D$l�D$(�D$t�D$ D�L$pD�D$D�T$@H�L$0�����H�|$x t!�D$ �   D�L$DD�D$@H�T$xH�L$0������V���3����]���H�D$8�L$d�HH�D$8�L$h�HH�D$8�L$H�HH�D$8�L$T�HH�D$8H�L$0H�H��$�   �@   �H��$�   �@    H���   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������H�T$H�L$H��   H�D$H����H��$�   ����H�D$ H��$�   �WL E3�A�   �?   H��������H�L$P����H�D$8H�D$8H�D$@L�D$@��  H�L$ �?����H�L$P�R���H��$�   �c���E3�A�   �?   H���I�����H�L$h�-���H�D$(H�D$(H�D$0L�D$0��  H�L$ ������H�L$h�����H�Ĉ   �������������������������������������������������������������������D�L$ L�D$H�T$H�L$H��8D�L$XL�D$PH�T$HH�L$@�m  �D$ �|$  u�D$ �gH�T$$H�L$P�J  ��u3��PH�D$@H�x tH�D$@H�H�z  ��v�  H�L$@H�A�|$$ tH�D$@H�PH�L$P��L  ��u3���D$ H��8���������������������������������������������������D�L$ D�D$H�T$H�L$H��8H�9� H�@0�L$`�L$ D�L$XD�D$PH�T$HH�L$@��   H��8�����������������������D�D$�T$H�L$H��(H�ߵ H�@ D�D$@�T$8H�L$0�PhH��(��������������D�L$ D�D$�T$H�L$H��8H��� H�@0�L$h�L$(�L$`�L$ D�L$XD�D$P�T$HH�L$@��  H��8���������������������������������L�D$�T$H�L$H��(H�/� H�@ L�D$@�T$8H�L$0�PpH��(��������������L�D$�T$H�L$H��(H�� H�@ L�D$@�T$8H�L$0���   H��(���������������������������L�D$H�T$H�L$H��HL�D$`H�T$XH�L$P�Yk  �D$0�|$0 u�D$0�pH�D$PH�x t
�D$4   ��D$4    �T$4H�L$`�<A  ��u3��<H�D$PH�x t,�D$    E3�A��� H�D$PH�PH�L$`�tC  ��u3���D$0H��H����������������������������������������������������D�L$ L�D$�T$H�L$H��8H�=��  ��   �D$X��t?H�|$@sH�D$    �
H�D$@H�D$ H��� H�@L�D$P�T$H�L$ ���  �P�=H�|$@sH�D$(   �
H�D$@H�D$(H�G� H�@L�D$P�T$H�L$(��P  ��D$X��H�L$@�  H��8�����������������H�L$H��8H�|$@ tMH�D$@H�D$ �=��  t(�   Hk��H�L$@�<�uH�D$@H��H����3 �H��� H�@H�L$ �H��8��������������H�L$H��(H�|$0 tH��� H�@H�L$0���  H��(���������������������H��(H�M� H�@�ﾭ����  H��(������������������H�L$H��(H�D$0H�8 tH�� H�@H�L$0H�	�H�D$0H�     H��(�������H�T$H�L$H��(H�ӱ H�@H�T$8H�L$0��X  H��(�������������������H�L$H�|$ t�   Hk��H�L$�<�u�   �3�����������������������H�T$H�L$H��(H�S� H�@H�T$8H�L$0��8  H��(�������������������H��(H�� H�@��@  H��(������̉T$H�L$H��8H�|$@s	H�D$@   H�D$@H��H����1 H�D$ H�|$  u3��G�|$H tH�D$@H��L��3�H�L$ �b� H�D$ � ����H�D$ H��H�D$ �A�    H�D$ H��8����H�L$H�D$H�     H�D$�@    H�D$H�@    H�D$�@    H�D$���������������������H�L$H��(H�L$0�  H��(���������H�L$H��xH�D$8����H�L$@�TQ  H�D$(H�D$(H�D$0H�T$0H��$�   �#   �D$ H�L$@�  �D$ H��x�������������H�T$H�L$H��XH�D$@����H�D$`H�x urL��� A�;   H��� �(   �����H�D$(H�|$( tH�T$hH�L$(�  H�D$0�	H�D$0    H�D$0H�D$8H�D$`H�L$8H�HH�D$`H�x u3��uH�D$`�x t#H�D$`H�8 t
�D$    ��D$     �D$ �GH�ޮ H�@xH�L$h�H�L$`H�H�D$`�@   H�D$`H�8 t
�D$$   ��D$$    �D$$H��X������������������H�L$H��8H�D$@�@   H�l� H�@x�PH�L$@H�H�D$@H�8 t
�D$    ��D$     �D$ H��8���������������̉T$H�L$H��(H�D$0H�8 uH�	� H�@(H� �H��� H�@x�T$8H�L$0H�	�PH��(����������H�L$H��(H�D$0�x t�   �/H�D$0H�x u3��H��� H�@xH�L$0H�QH�L$0H�	�P0H��(������������������H�L$H��HH�D$P�x t�   H�D$PH�8 t"H�M� H�@xH�L$PH�	�PH�D$PH�     H�D$PH�x tXH�D$PH�x t?H�D$PH�@H�D$(H�D$(H�D$ H�|$  t�   H�L$ �C  H�D$0�	H�D$0    H�D$PH�@    H��H�����������������̉L$H��(�T$0H�e� �x���H��(��������������������L�D$�T$H�L$H��   H�D$X�����D$4    ��$�   H�� �'���H��H�L$@�j����E3�H��� H�L$`�����E3�L�D$8H�T$`H�L$@�  ��u
�D$<   ��D$<    �D$<�D$0H�L$`�_����D$0��t,H��$�   ������D$4���D$4H�L$@�4���H��$�   �gA�   �T$8H�L$@�k  �D$ ����A�����L��$�   �T$8H�L$@��  H�T$@H��$�   �����D$4���D$4H�L$@�����H��$�   H�Ĉ   �����������������L�L$ L�D$�T$H�L$H��   H�D$x�����D$4    ��$�   H��� �����H��H�L$H�����E3�H�F� H�L$`�<����E3�L�D$8H�T$`H�L$H��  ��u
�D$<   ��D$<    �D$<�D$1H�L$`�
����D$1��t/H��$�   �w����D$4���D$4H�L$H�����H��$�   �2  A�   �T$8H�L$H�  �D$ ����A�����L��$�   �T$8H�L$H�  E3�H��� H��$�   �t����E3�L�D$8H��$�   H�L$H��  ��u
�D$@   ��D$@    �D$@�D$0H��$�   �<����D$0��t,H��$�   �����D$4���D$4H�L$H����H��$�   �gA�   �T$8H�L$H�H  �D$ ����A�����L��$�   �T$8H�L$H��  H�T$HH��$�   �r����D$4���D$4H�L$H����H��$�   H�Ĩ   ��������������L�L$ L�D$�T$H�L$H��   HǄ$�   �����D$0    ��$�   H��� ����H��H�L$H������E3�H�+� H�L$`�����E3�L�D$4H�T$`H�L$H�  ��u
�D$@   ��D$@    �D$@�D$:H�L$`������D$:��t/H��$�   �T����D$0���D$0H�L$H����H��$�   ��  A�   �T$4H�L$H��  �D$ ����A�����L��$�   �T$4H�L$H�l  E3�H�j� H�L$x�T����E3�L�D$4H�T$xH�L$H��  ��u
�D$<   ��D$<    �D$<�D$9H�L$x�"����D$9��t/H��$�   �����D$0���D$0H�L$H�����H��$�   �2  A�   �T$4H�L$H�+  �D$ ����A�����L��$�   �T$4H�L$H�  E3�H��� H��$�   �����E3�L�D$4H��$�   H�L$H�  ��u
�D$D   ��D$D    �D$D�D$8H��$�   �T����D$8��t,H��$�   ������D$0���D$0H�L$H�)���H��$�   �gA�   �T$4H�L$H�`
  �D$ ����A�����L��$�   �T$4H�L$H��  H�T$HH��$�   �����D$0���D$0H�L$H�����H��$�   H�ĸ   ����������������������L�L$ L�D$�T$H�L$H���   HǄ$�   �����D$4    ��$�   H��� ����H��H�L$@�����E3�H�G� H�L$h�)����E3�L�D$0H�T$hH�L$@�	  ��u
�D$\   ��D$\    �D$\�D$;H�L$h������D$;��t/H��$�   �d����D$4���D$4H�L$@�����H��$�   ��  A�   �T$0H�L$@� 	  �D$ ����A�����L��$�   �T$0H�L$@�|
  E3�H��� H��$�   �a����E3�L�D$0H��$�   H�L$@��  ��u
�D$X   ��D$X    �D$X�D$9H��$�   �)����D$9��t/H��$�   �����D$4���D$4H�L$@�����H��$�   �   A�   �T$0H�L$@�2  �D$ ����A�����L��$�   �T$0H�L$@�	  E3�H��� H��$�   �����E3�L�D$0H��$�   H�L$@�  ��u
�D$d   ��D$d    �D$d�D$:H��$�   �[����D$:��t/H��$�   ������D$4���D$4H�L$@�0���H��$�   �2  A�   �T$0H�L$@�d  �D$ ����A�����L��$   �T$0H�L$@��  E3�H��� H��$�   ������E3�L�D$0H��$�   H�L$@�N  ��u
�D$`   ��D$`    �D$`�D$8H��$�   �����D$8��t,H��$�   ������D$4���D$4H�L$@�b���H��$�   �gA�   �T$0H�L$@�  �D$ ����A�����L��$  �T$0H�L$@�  H�T$@H��$�   ������D$4���D$4H�L$@�����H��$�   H���   ���������������L�D$H�T$�L$H��8H�|$P tH�D$PH�D$ �H��� �  H�D$ L�D$ H�T$H�L$@�V� H��8������������������H�L$H��(H��� H�@xH�L$0�P H��(����������������H�T$H�L$H��HH�|$P u3��   H�T$PH�L$0�� �D$     H�D$(    L�D$(H�T$ H�L$0�� ��t]�|$ t�|$ u$H�L$(��  H�T$XH��������t�   �/�)�|$ u"H�L$(�x  H�T$XH���K  ��t�   ��3�H��H��������H�L$H���   HǄ$�   �����D$     E3�H�v� H��$�   �E���H�D$xH�D$xH�D$PH�L$P�����H�D$@H��$�   �)���H�|$@ u3��E  H�D$H    H�T$@H��$�   �t� L�D$8H�T$,H��$�   ��� ���  �|$,��   H�L$8��  H�D$0H�|$0 t~H��$�   �4���H�D$pH�D$pH�D$`�D$ ���D$ L�L$`A�   H��$�   H�L$0�  H�D$hH�D$hH�D$X�D$ ���D$ H��$�   H�L$X��  ��t
�D$(   ��D$(    �D$(�D$$�D$ ����t�d$ �H��$�   ������D$ ����t�d$ �H��$�   ������D$$��tH�D$8H�D$H������H�D$HH���   �������������������H�T$H�L$H���   HǄ$�   �����D$     H��$�    uWE3�H��� H��$�   �e���H�D$xH�D$xH�D$PH�L$P�����H��$�   H��$�   �F���H��$�    u3��  H�D$@    H��$�   H��$�   �� L�D$0H�T$(H��$�   �� ���A  �|$(��   H�L$0��  H�D$HH�|$H t~H��$�   �K���H�D$pH�D$pH�D$`�D$ ���D$ L�L$`A�   H��$�   H�L$H�  H�D$hH�D$hH�D$X�D$ ���D$ H��$�   H�L$X�
  ��t
�D$8   ��D$8    �D$8�D$$�D$ ����t�d$ �H��$�   �)�����D$ ����t�d$ �H��$�   �����D$$��tH�D$0H�D$@�@�9�|$(u2H�|$0 t*H�L$0�  H��$�   H���p   ��tH�D$0H�D$@�����H�D$@H���   ���������������H��(H�� H�@x�P(H��(����������H��(H��� ����H��(������������H�T$H�L$H��8H�T$HH�L$@�c   ��u
�D$    ��D$     �D$ H��8����̉T$H�L$H��(H�L$0�Y  �D$8����t
H�L$0�����H�D$0H��(�����������H�T$H�L$H��(H�S� H�@(H�T$8H�L$0���   H��(���D�D$�T$H�L$H��(H�� H�@(D�D$@�T$8H�L$0���   H��(�����������D�L$ L�D$H�T$H�L$H��(H�ٛ H�@(D�L$HL�D$@H�T$8H�L$0���   H��(���������������H�L$H�D$H� ���H�L$H��(H��� H��  H�L$0���   H��(����������L�L$ D�D$H�T$H�L$H��hH�D$8�����D$     H�8� H�@ L��$�   D��$�   H�T$@H�L$p��H  H�D$(H�D$(H�D$0H�T$0H�L$x�����D$ ���D$ H�L$@�T���H�D$xH��h����������������H�L$H��(H��� H��  H�L$0���   H��(����������D�L$ L�D$�T$H�L$H��8H�z� H�@(�L$`�L$ D�L$XL�D$P�T$HH�L$@���   H��8���������H�L$H�D$H�w� H�H�D$�������H�L$H�D$H�W� H�������������H�L$H��HH�D$PH�D$(H�|$( t@H�D$(H�D$0H�D$0H�D$ H�|$  tH�D$ H� �   H�L$ �H�D$8�	H�D$8    H�D$(    H��H��������H�L$H��(H��� H�@H�L$0��8  H��(�������������H�L$H��(H�X� H�@H�L$0��P  H��(�������������H�T$H�L$H��xH�D$8�����D$     H�� H�@H�T$@H��$�   ��@  H�D$(H�D$(H�D$0H�T$0H��$�   �2  �D$ ���D$ H�L$@�  H��$�   H��x�����������������H�L$H��(H��� H�@H�L$0��H  H��(������������̉T$�L$H��(H�e� H�@�T$8�L$0��(  H��(�������H�L$H��(H�8� H�@H�L$0��P  H��(�������������H��(H�� H�@��0  H��(�������D�D$�T$H�L$H��(H�ߗ H�@D�D$@�T$8H�L$0���  H��(�����������H�T$H�L$H��(H��� H�@H�T$8H�L$0���  H��(�������������������H�L$H��(H�h� H�@H�L$0���  H��(�������������H��(H�=� H�@���  H��(�������H�T$H�L$H��(H�� H�@H�T$8H�L$0���  H��(�������������������H�T$H�L$H��(H�Ӗ H�@H�T$8H�L$0���  H��(��̉T$H�L$H��(H�L$0�y����D$8����t
H�L$0�����H�D$0H��(�����������H��(H�m� H�@H���   H��(�������H�L$H��(H�H� H�@HH�L$0���   H��(�������������D�L$ L�D$H�T$H�L$H��(H�	� H�@HD�L$HL�D$@H�T$8H�L$0���   H��(���������������H�L$H��8H�D$ ����H�D$@H�������H��� H�@HH�L$@���   �H�D$@H��8����������������H�T$H�L$H��8H�D$ ����H�D$@H���Z����H�\� H�@HH�L$@���   H�F� H�@HH�T$HH�L$@���   �H�D$@H��8����������������H�T$H�L$H��8H�D$ ����H�D$@H��������H�� H�@HH�L$@���   H�֔ H�@HH�T$HH�L$@�P8�H�D$@H��8�������������������H�T$H�L$H��8H�D$ ����H�D$@H���z����H�|� H�@HH�L$@���   H�f� H�@HH�T$@H�L$H���   �H�D$@H��8����������������H�L$H��8H�D$ ����H�� H�@HH�L$@���   �H�D$@H���u���H��8����������������������H�T$H�L$H��(H�ӓ H�@HH�T$8H�L$0���   H��(�������������������L�L$ D�D$�T$H�L$H��8H��� H�@HH�L$`H�L$ L�L$XD�D$P�T$HH�L$@�P H��8����������H�L$H��(H�H� H�@HH�L$0�P(H��(����������������H�T$H�L$H��hH�D$8�����D$     H�� H�@HH�T$pH�L$@�P0H�D$(H�D$(H�D$0H�T$0H�L$x������D$ ���D$ H�L$@�1���H�D$xH��h�������������H�T$H�L$H��(H��� H�@HH�T$8H�L$0�P8H��(����������������������H�T$H�L$H��xH�D$8�����D$     H�B� H�@HH��$�   H�L$@�P@H�D$(H�D$(H�D$0H�T$0H��$�   �e����D$ ���D$ H�L$@�����H��$�   H��x��������������������H�T$H�L$H��xH�D$8�����D$     H��� H�@HH��$�   H�L$@�PHH�D$(H�D$(H�D$0H�T$0H��$�   ������D$ ���D$ H�L$@�0���H��$�   H��x��������������������H�T$H�L$H��xH�D$8�����D$     H�T$@H��$�   �?���H�D$(H�D$(H�D$0H��$�   H�L$0������D$ ���D$ H�L$@����H��$�   H��x�������������H�L$H��(H��� H�@HH�L$0�PPH��(����������������H�L$H��(H��� H�@HH�L$0���   H��(�������������H�T$H�L$H��(H�S� H�@HH�T$8H�L$0�PXH��(����������������������H�T$H�L$H��(H�� H�@HH�T$8H�L$0�P`H��(����������������������H�T$H�L$H��(H�ӏ H�@HH�T$8H�L$0�PhH��(����������������������H�T$H�L$H��(H��� H�@HH�T$8H�L$0�PpH��(����������������������D�D$H�T$H�L$H��(H�N� H�@HD�D$@H�T$8H�L$0���   H��(���������H�T$H�L$H��(H�� H�@HH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�ӎ H�@HH�T$8H�L$0���   H��(�������������������H�L$H��(H��� H�@HH�L$0���   H��(�������������H�T$H�L$H��(H�c� H�@HH�T$0H�L$8���   H�D$0H��(��������������L�D$H�T$H�L$H��hH�D$(�����D$     H�T$xH�L$0�]����H��� H�@HH��$�   H�L$0���   H�T$0H�L$p�/����D$ ���D$ H�L$0����H�D$pH��h�����������������H�T$H�L$H��(H��� H�@HH�T$8H�L$0���   H�D$0H��(��������������H�T$H�L$H��(H�S� H�@HH�T$8H�L$0�PxH��(����������������������H�T$H�L$H��8H�� H�@HH�T$HH�L$@�Px��u
�D$    ��D$     �D$ H��8������������H�T$H�L$H��hH�D$8�����D$     H��� H�@HH�T$pH�L$@���   H�D$(H�D$(H�D$0H�T$0H�L$x訹���D$ ���D$ H�L$@�޹��H�D$xH��h����������D�L$ D�D$H�T$H�L$H��HH�9� H�@P��$�   �L$0�L$x�L$(�L$p�L$ D�L$hD�D$`H�T$XH�L$P�P H��H�������H�L$H��(H�� H�@PH�L$0�P(H��(���������������̉T$H�L$H��(H��� H�@P�T$8H�L$0�P0H��(��������D�L$ D�D$H�T$H�L$H��(H�y� H�@PD�L$HD�D$@H�T$8H�L$0�P8H��(������������������D�D$H�T$H�L$H��(H�.� H�@PD�D$@H�T$8H�L$0�P@H��(������������D�D$H�T$H�L$H��(H�� H�@PA�   D�D$@H�T$8H�L$0�P8H��(����������������������D�D$H�T$H�L$H��(H��� H�@PD�D$@H�T$8H�L$0�PHH��(������������H�L$H��(H�h� H�@PH�L$0�PPH��(����������������H�L$H��(H�8� H�@PH�L$0�PXH��(����������������H�L$H��(H�� H�@PH�L$0�P`H��(���������������̉T$H�L$H��(H�ԉ H�@P�T$8H�L$0�PhH��(��������H�T$H�L$H��(H��� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�c� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�#� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�c� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�#� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�c� H�@PH�T$8H�L$0��  H��(�������������������H�T$H�L$H��XH�D$(����H�L$0�����H�T$0H�L$`�   ��u�D$     H�L$0�d����D$ �%H�T$0H�L$h�4����D$$   H�L$0�=����D$$H��X����������H�T$H�L$H��8H�T$ H�L$@�������u3��+�D$ ��t
�D$$   ��D$$    H�D$H�L$$��   H��8������������H�T$H�L$H��hH�D$@�����D$     H�D$(    H�T$ H�L$p�i�����u3���   �|$  u=H�L$H�����H�D$0H�D$0H�D$8H�T$8H�L$x�*  �H�L$H�O����   �   H�˅ H�@L�0� �j  �L$ ���  H�D$(H�|$( u�����H�L$p����3��SE3�D�D$ H�T$(H�L$p�������uH�L$(�D���3��*�D$ ��E3�D��H�T$(H�L$x�*  H�L$(�����   H��h������������������H�T$H�L$H��8H�D$HH��H�L$@�������t>H�D$HH��H��H�L$@������t$H�D$HH��H��H�L$@������t
�D$    ��D$     �D$ H��8��������������H�T$H�L$H��8H�D$HH��H�L$@������t>H�D$HH��H��H�L$@�v�����t$H�D$HH��H��H�L$@�\�����t
�D$    ��D$     �D$ H��8��������������H�T$H�L$H��8H�D$HH��H�L$@�������tXH�D$HH��H��H�L$@�������t>H�D$HH��H��H�L$@������t$H�D$HH��$H��H�L$@������t
�D$    ��D$     �D$ H��8��������������������H�T$H�L$H��8H�D$HH��H�L$@�������tXH�D$HH��H��H�L$@������t>H�D$HH��0H��H�L$@������t$H�D$HH��HH��H�L$@�r�����t
�D$    ��D$     �D$ H��8�������������������̈T$H�L$H��(H�Ԃ H�@P�T$8H�L$0�PpH��(������̈T$H�L$H��(H��� H�@P�T$8H�L$0�PxH��(�������f�T$H�L$H��(H�s� H�@P�T$8H�L$0���   H��(�������������������f�T$H�L$H��(H�3� H�@P�T$8H�L$0���   H��(������������������̉T$H�L$H��(H�� H�@P�T$8H�L$0���   H��(��������������������̉T$H�L$H��(H��� H�@P�T$8H�L$0���   H��(����������������������L$H�L$H��(H�r� H�@P�L$8H�L$0���   H��(������������������L$H�L$H��(H�2� H�@P�L$8H�L$0���   H��(�����������������H�T$H�L$H��(H�� H�@PH�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��� H�@PH�T$8H�L$0��  H��(�������������������H�T$H�L$H��hH�D$8����H�T$@H�L$x�:���H�D$(H�D$(H�D$0H�T$0H�L$p�l   �D$ H�L$@詭���D$ H��h���������������������̉T$H�L$H��8�|$H t�D$ ��D$  �T$ H�L$@����H��8�������������H�T$H�L$H��H3�H�L$X��$  ���D$ H�� H�@L�>� ��  �L$ ���  H�D$0H�|$0 u�����H�L$P����3��iE3�D�D$ H�T$0H�L$X�H$  �T$ H�L$P�J�����t"D�D$ H�T$0H�L$P�������t
�D$$   ��D$$    �D$$�D$(H�L$0������D$(H��H������������������H�T$H�L$H��8H�D$H�H�L$@�O�����t:H�D$H�HH�L$@�7�����t"H�D$H�HH�L$@������t
�D$    ��D$     �D$ H��8�����������������H�T$H�L$H��8H�D$H�H�L$@������t:H�D$H�HH�L$@�������t"H�D$H�HH�L$@�������t
�D$    ��D$     �D$ H��8�����������������H�T$H�L$H��8H�D$HH��H�L$@�������tXH�D$HH��H��H�L$@�������t>H�D$HH��H��H�L$@������t$H�D$HH��$H��H�L$@������t
�D$    ��D$     �D$ H��8��������������������H�T$H�L$H��8H�D$HH��H�L$@�������tXH�D$HH��H��H�L$@������t>H�D$HH��0H��H�L$@������t$H�D$HH��HH��H�L$@�r�����t
�D$    ��D$     �D$ H��8��������������������H��(H��| H�@P�H��(�����������H�L$H��(H��| H�@PH�L$0H�	�PH�D$0H�     H��(�����������������D�L$ L�D$H�T$H�L$H��hH�9| H�@P��$�   �L$P��$�   �L$H��$�   �L$@��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ D��$�   L��$�   H�T$xH�L$p��   H��h������������D�L$ L�D$H�T$H�L$H��8H��{ H�@P�L$`�L$ D�L$XL�D$PH�T$HH�L$@�PH��8����������H��(H�]{ H�@P�PH��(����������H�L$H��(H�8{ H�@PH�L$0H�	�PH�D$0H�     H��(�����������������D�D$H�T$H�L$H��(H��z H�@XD�D$@H�T$8H�L$0�PH��(������������H�L$H��(H��z H�@XH�L$0�PH��(����������������H�L$H��(H��z H�@XH�L$0�P0H��(����������������H�L$H��(H�Xz H�@XH�L$0�P(H��(����������������H�L$H��(H�(z H�@XH�L$0�P@H��(����������������H�L$H��(H��y H�@XH�L$0�PPH��(����������������H�L$H��(H��y H�@XH�L$0�PHH��(����������������L�D$�T$H�L$H��(H��y H�@XL�D$@�T$8H�L$0�P8H��(��������������H�T$H�L$H��xH�D$8�����D$     H�By H�@XH�T$@H��$�   �P H�D$(H�D$(H�D$0H�T$0H��$�   �e����D$ ���D$ H�L$@�����H��$�   H��x��������������������H��(H��x H�@X3�3��H��(�������H�L$H��(H��x H�@XH�L$0H�	�PH�D$0H�     H��(�����������������H�L$H��(H�hx H�@XH�L$0�PhH��(����������������H�L$H��(H�8x H�@XH�L$0�PpH��(����������������H�T$H�L$H��xH�D$8�����D$     H��w H�@XH�T$@H��$�   �PxH�D$(H�D$(H�D$0H�T$0H��$�   �����D$ ���D$ H�L$@�p���H��$�   H��x��������������������L�D$H�T$H�L$H��hH�D$8�����D$     H�]w H�@XL��$�   H�T$@H�L$p���   H�D$(H�D$(H�D$0H�T$0H�L$x�K����D$ ���D$ H�L$@聤��H�D$xH��h�������������H��(H��v H�@X�PXH��(����������H�L$H��(H��v H�@XH�L$0H�	�P`H�D$0H�     H��(�����������������L�D$H�T$H�L$H��(H�~v H�@L�D$@H�T$8H�L$0��  H��(���������L�D$H�T$H�L$H��(H�>v H�@L�D$@H�T$8H�L$0��  H��(���������L�D$H�T$H�L$H��(H��u H�@L�D$@H�T$8H�L$0��  H��(���������L�D$H�T$H�L$H��(H��u H�@L�D$@H�T$8H�L$0��   H��(��������̈T$H�L$H��(H��u H�@�T$8H�L$0�PH��(������̈T$H�L$H��(H�Tu H�@�T$8H�L$0�PH��(�������f�T$H�L$H��(H�#u H�@�T$8H�L$0�P H��(����������������������f�T$H�L$H��(H��t H�@�T$8H�L$0�P(H��(���������������������̉T$H�L$H��(H��t H�@�T$8H�L$0�P0H��(�������̉T$H�L$H��(H�tt H�@�T$8H�L$0�P8H��(��������H�T$H�L$H��(H�Ct H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�t H�@H�T$8H�L$0��   H��(��������������������L$H�L$H��(H��s H�@�L$8H�L$0�P@H��(���������������������L$H�L$H��(H��s H�@�L$8H�L$0�PHH��(���������������������L$H�L$H��(H�Bs H�@�L$8H�L$0�PPH��(�������������������̉T$H�L$H��(H�s H�@�T$8H�L$0�PXH��(��������H�T$H�L$H��(H��r H�@H�T$8H�L$0�P`H��(����������������������H�T$H�L$H��(H��r H�@H�T$8H�L$0�PhH��(����������������������H�T$H�L$H��(H�Sr H�@H�T$8H�L$0�PpH��(����������������������H�T$H�L$H��(H�r H�@H�T$8H�L$0�PxH��(����������������������H�T$H�L$H��(H��q H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��q H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�Sq H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�q H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��p H�@H�T$8H�L$0���   H��(�������������������L�L$ D�D$H�T$H�L$H��8H��p H�@�L$`�L$ L�L$XD�D$PH�T$HH�L$@���  H��8�������H�T$H�L$H��(H�Cp H�@H�T$8H�L$0��  H��(�������������������H�T$H�L$H��(H�p H�@H�T$8H�L$0���   H��(�������������������D�D$H�T$H�L$H��(H��o H�@D�D$@H�T$8H�L$0���   H��(���������H�T$H�L$H��(H�|$8 u3��H�wo H�@@H�T$8H�L$0�PP�   H��(���������������������D�L$ D�D$H�T$H�L$H��8H�)o H�@�L$`�L$ D�L$XD�D$PH�T$HH�L$@���  H��8�������H�T$H�L$H��(H��n H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��n H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�cn H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�#n H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��m H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��m H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�cm H�@H�T$8H�L$0��p  H��(�������������������H�T$H�L$H��(H�#m H�@H�T$8H�L$0��  H��(�������������������H�T$H�L$H��(H��l H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H��l H�@H�T$8H�L$0���   H��(�������������������H�T$H�L$H��(H�cl H�@H�T$8H�L$0��   H��(�������������������H�T$H�L$H��(H�#l H�@H�T$8H�L$0��  H��(�������������������H�T$H�L$H��(H��k H�@H�T$8H�L$0��  H��(�������������������H�T$H�L$H��(H��k H�@H�T$8H�L$0��  H��(�������������������H�T$H�L$H��(H�ck H�@H�T$8H�L$0��   H��(�������������������H�T$H�L$H��(H�#k H�@H�T$8H�L$0��(  H��(�������������������H�T$H�L$H��(H��j H�@H�T$8H�L$0��0  H��(�������������������H�T$H�L$H��(H��j H�@H�T$8H�L$0��8  H��(�������������������H�T$H�L$H��(H�cj H�@H�T$8H�L$0��@  H��(�������������������H�T$H�L$H��(H�#j H�@H�T$8H�L$0��H  H��(�������������������H�T$H�L$H��(H��i H�@H�T$8H�L$0��P  H��(�������������������H�T$H�L$H��(H��i H�@H�T$8H�L$0��X  H��(�������������������H�T$H�L$H��(H�ci H�@H�T$8H�L$0��  H��(�������������������D�D$H�T$H�L$H��(H�i H�@D�D$@H�T$8H�L$0��`  H��(���������L�D$H�T$H�L$H��(H��h H�@L�D$@H�T$8H�L$0��h  H��(���������H�T$H�L$H��8H�|$H t&H��h H�@@H�T$HH�L$@�PH��t
�D$    ��D$     �D$ H��8��������������������D�D$H�T$H�L$H��(H�>h H�@@L�D$0�T$@H�L$8���   H��(����������D�L$ D�D$H�T$H�L$H��8H��g H�@�L$`�L$ D�L$XD�D$PH�T$HH�L$@���  H��8�������H�L$H��(H��g H�@H�L$0��x  H��(������������̉T$H�L$H��(H��g H�@�T$8H�L$0���  H��(���������������������H�T$H�L$H��(H�Cg H�@H�T$8H�L$0���  H��(������������������̉T$H�L$H��(H�g H�@�T$8H�L$0���  H��(���������������������D�D$�T$H�L$H��(H��f H�@D�D$@�T$8H�L$0���  H��(�����������H�L$H��(H��f H�@H�L$0���  H��(�������������L�D$H�T$H�L$H��(H�Nf H�@L�D$@H�T$8H�L$0���  H��(���������H�L$H��(H�f H�@H�L$0���  H��(�������������H�L$H��(H��e H�@H�L$0���  H��(�������������H�L$H��(H��e H�@H�L$0���  H��(�������������H�L$H��(H��e H�@H�L$0���  H��(�������������H��(H�]e H�@���  H��(�������H�L$H��(H�8e H�@H�L$0���  H�D$0H�     H��(�����������������D�L$ L�D$�T$H�L$H��8H��d H�@�L$`�L$ D�L$XL�D$P�T$HH�L$@�H��8�������������H�L$H��(H��d H�@H�L$0�PH��(����������������D�L$ L�D$H�T$H�L$H��8H�id H�@H�L$`H�L$ D�L$XL�D$PH�T$HH�L$@���  H��8���������������������D�L$ L�D$H�T$H�L$H��(H�	d H�@D�L$HL�D$@H�T$8H�L$0��   H��(��������������̉T$H�L$H��(H��c H�@�T$8H�L$0�PH��(��������L�D$H�T$H�L$H��(H��c H�@L�D$@H�T$8H�L$0�PH��(�����������̉T$H�L$H��(H�Tc H�@�T$8H�L$0�P H��(��������D�D$H�T$H�L$H��(H�c H�@D�D$@H�T$8H�L$0�P(H��(������������H�T$H�L$H��(H��b H�@H�T$8H�L$0�P0H��(����������������������H�T$H�L$H��(H��b H�@H�T$8H�L$0���  H��(�������������������H�L$H��(H�hb H�@H�L$0�P8H��(����������������H�L$H��hH�D$0����H�T$8H�L$p�����H�L$8�������u�D$     H�L$8������D$ �   �   H�L$8������u&H�L$8������u�D$$    H�L$8�����D$$�O�   H�L$p�������u&H�L$p�/�����u�D$(    H�L$8�Y����D$(��D$,   H�L$8�A����D$,H��h���������H�L$H��(H�Xa H�@H�L$0�P@H��(����������������H�T$H�L$H��(H�#a H�@H�T$8H�L$0�PPH��(����������������������L�L$ D�D$H�T$H�L$H��8H��` H�@H�L$`H�L$ L�L$XD�D$PH�T$HH�L$@��   H��8���������������������L�L$ L�D$H�T$H�L$H��(H�y` H�@L�L$HL�D$@H�T$8H�L$0��   H��(���������������H�L$H��(H�8` H�@H�L$0��  H��(�������������D�D$�T$H�L$H��(H��_ H�@D�D$@�T$8H�L$0��  H��(�����������H�L$H��xH�D$8�����D$     H��_ H�@H�L$@�PHH�D$(H�D$(H�D$0H�T$0H��$�   ������D$ ���D$ H�L$@�=���H��$�   H��x�����������������H�L$H��xH�D$8�����D$     H�7_ H�@H�L$@���  H�D$(H�D$(H�D$0H�T$0H��$�   �_����D$ ���D$ H�L$@����H��$�   H��x��������������H�L$H��8�D$     �   H�L$@�0  �D$ ���D$ H�D$@H��8������������H�L$H��   H�D$X�����D$     H�=�^  t:H��$�   H�z^ �����H�D$PH�D$PH�D$@�D$ ���D$ H�D$@H�D$(�.H�L$`�U���H�D$0H�D$0H�D$H�D$ ���D$ H�D$HH�D$(H�D$(H�D$8H�T$8H��$�   �E����D$ ���D$ �D$ ����t�d$ �H�L$`������D$ ����t�d$ �H��$�   �r���H��$�   H�ĸ   ������������������̉T$H�L$H��xH�D$8�����D$     H�c] H�@��$�   H�L$@���  H�D$(H�D$(H�D$0H�T$0H��$�   �����D$ ���D$ H�L$@�����H��$�   H��x�������������������L�D$�T$H�L$H��(H��\ H�@L�D$@�T$8H�L$0���  H��(�����������L�D$�T$H�L$H��(H��\ H�@L�D$@�T$8H�L$0���  H��(�����������H�L$H��(H�h\ H�@H�L$0���  H��(�������������D�D$H�T$H�L$H��hH�D$8�����D$     H�\ H�@D��$�   H�T$xH�L$@���  H�D$(H�D$(H�D$0H�T$0H�L$p�����D$ ���D$ H�L$@�A���H�D$pH��h������������̉T$H�L$H��(H��[ H�@�T$8H�L$0���  H��(���������������������H�T$H�L$H��(H�c[ H�@H�T$8H�L$0���  H��(���H�T$H�L$H��(H�3[ H�@(H�T$0H�L$8�P8H�D$0H��(�D�L$ D�D$H�T$H�L$H��(H��Z H�@(D�L$HD�D$@H�T$8H�L$0���   H��(��������������̉T$H�L$H��(H��Z H�@(�T$8H�L$0���   H��(�����D�L$ D�D$H�T$H�L$H��(H�yZ H�@(D�L$HD�D$@H�T$8H�L$0�P H��(��H�L$H�D$H�@    H�D$�     H�D$�@    H�D$�@   H�D$����������������������D�L$ D�D$H�T$H�L$H��(H��Y H���   D�L$HD�D$@H�T$8H�L$0�P(H��(���������������H�T$H�L$H��(H��Y H���   H�T$8H�L$0�P0H��(�������������������D�D$H�T$H�L$H��(H�^Y H���   D�D$@H�T$8H�L$0�P8H��(���������H�T$H�L$H��(H�#Y H���   H�T$8H�L$0�P@H��(�������������������D�D$H�T$H�L$H��(H��X H��  D�D$@H�T$8H�L$0�P0H��(���������D�L$ L�D$H�T$H�L$H��(H��X H��  D�L$HL�D$@H�T$8H�L$0�P8H��(���������������D�L$ L�D$H�T$H�L$H��(H�IX H��  D�L$HL�D$@H�T$8H�L$0�P@H��(���������������H�L$H��(H�X H��  H�L$0�PHH��(�������������D�L$ L�D$H�T$H�L$H��8H��W H��  H�L$`H�L$ D�L$XL�D$PH�T$HH�L$@���  H��8������������������L�L$ L�D$H�T$H�L$H��(H�iW H��  L�L$HL�D$@H�T$8H�L$0���  H��(������������H�T$H�L$H��(H�#W H���   H�T$8H�L$0���   H��(����������������H�L$H��(H��V H���   H�L$0���   H��(���������̉T$H�L$H��(H��V H��  �T$8H�L$0���  H��(������������������D�D$�T$H�L$H��(H�oV H��  D�D$@�T$8H�L$0���  H��(��������H�L$H��(H�8V H���   H�L$0��P  H��(����������L�L$ L�D$H�T$H�L$H��(H�|$8 u�AH�|$H tH�T$HH�L$8�  �(H�|$@ tH�T$@H�L$8�  �H�T$0H�L$8�  H��(���������H��(H��U H���   �P`H��(�������H�L$H��(H�D$0H�8 tH�mU H���   H�L$0H�	�P H�D$0H�     H��(������������������̉T$H�L$H��8H�$U H���   H�L$@�P�D$ �D$H�L$ #ȋ���t�D$H�ЋL$ #ȋ��D$ ��D$H�L$ ȋ��D$ H��T H���   �T$ H�L$@�PH��8�������L�L$ L�D$H�T$H�L$H��HH��T H��  ��$�   �L$0�D$x�D$(H�L$pH�L$ L�L$hL�D$`H�T$XH�L$P���  H��H�����������L�L$ L�D$H�T$H�L$H��8H�)T H��  �L$h�L$(H�L$`H�L$ L�L$XL�D$PH�T$HH�L$@��   H��8����������H�L$H��(H��S H���   H�L$0��X  H��(����������H�T$H�L$H��(H��S H���   H�T$8H�L$0���  H��(����������������H�L$H��(H�hS H���   H�L$0���   H��(����������H�T$H�L$H��(H�3S H���   H�T$8H�L$0���   H��(����������������D�D$H�T$H�L$H��(H��R H���   D�D$@H�T$8H�L$0���   H��(����������������������H�L$H��(H��R H���   H�L$0���   H��(����������H�T$H�L$H��(H�sR H���   H�T$8H�L$0���   H��(����������������H�T$H�L$H��(H�3R H���   H�T$8H�L$0���   H��(����������������D�D$H�T$H�L$H��(H��Q H���   D�D$@H�T$8H�L$0���   H��(����������������������L�D$H�T$H�L$H��(H��Q H���   L�D$@H�T$8H�L$0��P  H��(����������������������H�L$H��(H�XQ H���   H�L$0���   H��(����������H�L$H��(H�(Q H���   H�L$0���   H��(����������H�T$H�L$H��(H��P H���   H�T$8H�L$0���   H��(����������������H�L$H��(H��P H���   H�L$0��  H��(����������H�T$H�L$H��(H��P H���   H�T$8H�L$0��   H��(����������������H�L$H��(H�HP H���   H�L$0��   H��(����������H�L$H��(H�P H��  H�L$0���   H��(����������H�T$H�L$H��(H��O H���   H�T$8H�L$0��  H��(����������������D�L$ D�D$H�T$H�L$H��8H��O H���   H�L$`H�L$ D�L$XD�D$PH�T$HH�L$@��(  H��8������������������D�L$ L�D$H�T$H�L$H��(H�9O H���   D�L$HL�D$@H�T$8H�L$0��0  H��(������������D�L$ L�D$H�T$H�L$H��(H��N H���   D�L$HL�D$@H�T$8H�L$0��8  H��(������������D�D$H�T$H�L$H��(H��N H���   D�D$@H�T$8H�L$0��@  H��(����������������������D�D$H�T$H�L$H��(H�NN H���   D�D$@H�T$8H�L$0��H  H��(���������������������̉L$H��(H�	N H���   �L$0��  H��(������������H�L$H��(H�D$0H�8 tH��M H���   H�L$0H�	�P H�D$0H�     H��(�������������������H��(H��M H���   �P`H��(������̉L$H��(H�iM H���   A�   H�T$03��PhH��(���������������������̉L$H��(H�)M H���   A�   H�T$0�   @�PhH��(������������������̉T$H�L$H��(H��L H���   D�D$8H�T$03��PhH��(������������������H��(H��L H���   �H��(��������H�L$H��(H�D$0H�8 tH�}L H���   H�L$0H�	�PH�D$0H�     H��(�������������������H��(H�=L H���   �P@H��(�������H�L$H��(H�D$0H�8 tH�L H���   H�L$0H�	�PPH�D$0H�     H��(�������������������L�L$ D�D$H�T$H�L$H��(H��K H�@@L�L$HD�D$@H�T$8H�L$0���   H��(���������������L�L$ D�D$�T$H�L$H��8�|$PqF t�>H�D$XH�D$ H�|$  u�*H�T$@H�L$ �*  H�L$@�x��L�D$ �T$HH���O  H��8�����������H�T$H�L$H��(H�K H�@H�T$8H�L$0���  H��(�������������������H�T$H�L$H��8H�L$H�x��A����E  H����z H�D$ H�L$@��w��A����E  H���z H��J H�IH�L$(H�T$ H��H�D$(���  H��8������������H�T$H�L$H��(H�CJ H��  H�T$8H�L$0���   H��(����������������H�T$H�L$H��(H�J H��  H�T$8H�L$0���   H��(����������������L�D$�T$H�L$H��(H��I H�@ L�D$@�T$8H�L$0���   H��(�����������H�T$H�L$�   �����������������H�T$H�L$����������������������D�L$ L�D$H�T$H�L$�   �������L�D$H�T$H�L$�   ������������L�L$ D�D$H�T$H�L$�   �������L�L$ L�D$H�T$H�L$�   �������L�D$H�T$H�L$�����������������H�T$H�L$3���������������������D�L$ L�D$H�T$H�L$3�����������D�D$H�T$H�L$3����������������L�L$ L�D$H�T$H�L$3�����������L�L$ L�D$H�T$H�L$�   �������L�L$ L�D$H�T$H�L$�   �������L�L$ L�D$H�T$H�L$�   �������L�L$ L�D$H�T$H�L$3�����������L�D$H�T$H�L$3����������������L�L$ L�D$�T$H�L$H�D$H�L$H�HhH�D$H�c���H�HH�D$H�/  H�HpH�D$H�'  H�HxH�D$H�  H���   H�D$H�  H���   H�D$H�  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$H��  H���   H�D$�L$(�H@H�D$�L$�H�D$H�L$ H�H`H�D$H�L$0H�HPH�D$H�@X    ���������������������L�L$ D�D$H�T$�L$H��x  E3��@  H�L$0�  H�D$(    ��$�  �D$ L��$�  L��$�  ��$�  H�L$0�����H��$�  H��$�   �D$ @  L�L$0L��$�  ��$�  �   �� H��x  ������������������H�T$H�L$H��X  H�D$h������  H��$`  H�H��$`  H�8 u�a  H��$h  H��$�   �ί���E3�H�3� H�L$p�5r��H�D$PH�D$PH�D$`H�T$`H��$�   蘯���H��$(  �
���H�D$XH�D$XH�D$HL��$�   H�T$HH��$   �A���H�D$8H�D$8H�D$@L��$�   H�T$@H��$�   ����H�D$(H�D$(H�D$0E3�A�����H�T$0H��$`  H��	  ��t
�D$$   ��D$$    �D$$�D$ H��$�   辯���H��$   谯���H��$(  袯���H��$�   蔯���H�L$p�4q���H��$�   �{����D$ ��tH��$`  H���r  H��$`  H��X  ������������������̉T$H�L$H��(�L$8��   H�L$0H�H�D$0H��(���������H�L$H��(H�D$0H���
  H��(��H��`��H��`��H��`��H��` ��H��`(��H��`0��H��`8��H��`@��H��`H��H��`P��H��`X��H��``��H��`h��H��`p��H��`x��H����   ���D�D$�T$H�L$H��(HcD$8�L$@���   L����H�L$0�2H H��(������������H��(H�]B H�@0��@  H��(�������H�L$H��(H�8B H�@0H�L$0H�	��H  H�D$0H�     H��(��������������H�T$H�L$H��(H��A H�@0H�T$0H�L$8��P  H�D$0H��(��������������H�T$H�L$H��(H��A H�@0H�T$0H�L$8��X  H��(�������������������H�T$H�L$H��8H�sA H�@0H�T$@H�L$H��X  ��u
�D$    ��D$     �D$ H��8���������H�T$H�L$H��8H�|$H tH�L$H�p&  H�D$ �	H�D$     H�A H�@0H�T$ H�L$@��p  H��8�����������������H�T$H�L$H��(H��@ H�@0H�T$8H�L$0��x  H��(�������������������L�D$H�T$H�L$H��(H�~@ H�@0L�D$@H�T$8H�L$0���  H��(���������L�D$H�T$H�L$H��(H�>@ H�@0L�D$@H�T$8H�L$0���  H��(���������H�T$H�L$H��(H�@ H�@0H�T$8H�L$0���  H��(�������������������D�D$H�T$H�L$H��hH�D$8�����D$     H��? H�@0D��$�   H�T$pH�L$@���  H�D$(H�D$(H�D$0H�T$0H�L$x�l���D$ ���D$ H�L$@��l��H�D$xH��h�������������H�L$H��(H�8? H�@0H�L$0���  H��(�������������H�L$H��(H�? H�@0H�L$0���  H��(������������̉T$H�L$H��(H��> H�@0�T$8H�L$0���  H��(��������������������̉T$H�L$H��(H��> H�@0�T$8H�L$0���  H��(���������������������H��(H�]> H�@0��`  H��(�������H��(H�=> H�@0��h  H��(�������H��(H�> H�@0���  H��(�������H��(H��= H�@0���  H��(�������H��(H��= H�@0���  H��(�������H�L$H��(H��= H�@0H�L$0H�	���  H�D$0H�     H��(��������������D�L$ L�D$�T$H�L$H��8H�j= H�@0�L$h�L$(H�L$`H�L$ D�L$XL�D$P�T$HH�L$@���  H��8���������������D�L$ L�D$H�T$H�L$H��8H�	= H�@0�L$h�L$(�L$`�L$ D�L$XL�D$PH�T$HH�L$@���  H��8���������������H�L$H��(H��< H�@0H�L$0�PH��(����������������D�L$ D�D$�T$H�L$H��8H�z< H�@0�L$`�L$ D�L$XD�D$P�T$HH�L$@���   H��8���������H�T$H�L$H��(H�3< H�@0H�T$8H�L$0���   H��(�������������������H�L$H��(H��; H�@0H�L$0�P@H��(����������������H�L$H��XH�D$8����H��; H�@0A��  H�T$`H�L$@��X  H�D$(H�D$(H�D$0H�L$0�D!  �D$ H�L$@�F  �D$ H��X��������������L�L$ D�D$H�T$H�L$H��8H�I; H�@0H�L$`H�L$ L�L$XD�D$PH�T$HH�L$@��   H��8���������������������L�L$ D�D$H�T$H�L$H��(H��: H�@0L�L$HD�D$@H�T$8H�L$0�P8H��(������������������D�L$ D�D$�T$H�L$H��8H��: H�@0�L$`�L$ D�L$XD�D$P�T$HH�L$@���  H��8���������L�L$ D�D$H�T$H�L$H��8H�I: H�@0�L$`�L$ L�L$XD�D$PH�T$HH�L$@�PHH��8����������D�L$ D�D$�T$H�L$H��8H��9 H�@0�L$`�L$ D�L$XD�D$P�T$HH�L$@�PPH��8������������D�L$ D�D$H�T$H�L$H��8H��9 H�@0�L$`�L$ D�L$XD�D$PH�T$HH�L$@�PXH��8����������D�L$ D�D$H�T$H�L$H��XH�Y9 H�@0��$�   �L$H��$�   �L$@��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ D�L$xD�D$pH�T$hH�L$`���   H��X�������������D�L$ D�D$�T$H�L$H��XH�L$`�e���ȉD$@H�L$`��e����H��8 H�I0H�L$H�T$x�T$8�T$p�T$0�T$h�T$(�T$@�T$ D��E3�3�H�L$`H�D$H�PhH��X��������������������D�L$ D�D$�T$H�L$H��HH�:8 H�@0��$�   �L$8��$�   �L$0�L$x�L$(�L$p�L$ D�L$hD�D$`�T$XH�L$P�PhH��H��������������D�D$�T$H�L$H��(H��7 H�@0D�D$@�T$8H�L$0���   H��(�����������H�T$H�L$H��(H��7 H�@0H�T$8H�L$0���   H��(�������������������H�L$H��(H�X7 H�@0H�L$0���   H��(�������������H�L$H��(H�(7 H�@0H�L$0���   H��(�������������H�L$H��(H��6 H�@0H�L$0���   H��(������������̉T$H�L$H��(H��6 H�@0�T$8H�L$0���   H��(��������������������̉T$H�L$H��(H��6 H�@0�T$8H�L$0���   H��(���������������������H�L$H��(H�H6 H�@0H�L$0���   H��(�������������L�D$�T$H�L$H��(H�6 H�@0L�D$@�T$8H�L$0���  H��(�����������L�L$ D�D$H�T$H�L$H��XH�D$8�����D$     H��5 H�@0L�L$xD�D$pH�T$`H�L$@��x  H�D$(H�D$(H�D$0H�T$0H�L$h�D  �D$ ���D$ H�L$@�/  H�D$hH��X����������������������H��(H�=5 H�@0�H��(�����������H�L$H��(H�5 H�@0H�L$0H�	�PH�D$0H�     H��(�����������������D�L$ D�D$H�T$H�L$H��8H��4 H�@0�L$h�L$(�L$`�L$ D�L$XD�D$PH�T$HH�L$@���  H��8���������������H�L$H��(H�x4 H�@0H�L$0H�	�PH�D$0H�     H��(�����������������D�D$H�T$H�L$H��8H�L$H��  H�L$@�������uH�Ƅ ��  �t  3��   H�D$(    H��3 H�@0L�L$$L�D$(�T$PH�L$@���  ��u3��]�D$     �
�D$ ���D$ �D$$9D$ }0HcD$ H�L$(H�<� u��HcD$ H�L$(H��H��H�L$H��  �H�L$(�P����   H��8�������D�D$H�T$H�L$H��HH�L$X�S  H�L$P�������uH�� ��  �  3��   H�D$(    H�3 H�@0L�L$$L�D$(�T$`H�L$P���  ��u3��   H�|$( u3��{�D$     �
�D$ ���D$ �D$$9D$ }NHcD$ H�L$(H�<� tHcD$ H�L$(H���G�����u��HcD$ H�L$(H��H�D$0H�T$0H�L$X�?  �H�L$(�C����   H��H����������D�D$H�T$H�L$H��(H�>2 H�@0D�D$@H�T$8H�L$0���  H��(���������H�L$H��(H�2 H�@0H�L$0���  H��(�������������H�L$H��(H��1 H�@0H�L$0���  H��(�������������H�T$H�L$H��(H��1 H�@0H�T$8H�L$0���  H��(�������������������H��(H�m1 H�@0���  H��(�������H�L$H��(H�H1 H�@0H�L$0H�	���  H�D$0H�     H��(��������������H�L$H��8H�D$ ����H�D$@H��H���m  �H�L$@�R   �H�D$@H��8��������H�L$H��8H�D$ ����H�L$@�   �H�D$@H��H���R  H��8��������������H�L$H�D$H�     H�D$Hǀ�       H�D$ǀ�       H�D$ǀ�       H�D$W����   H�D$ǀ�   ����H�D$ǀ�      �������������������H�L$H��8H�D$@H�8 t6H�D$@H���D$     E3�A�   H��H�D$@H��"  H�D$@H�     H�D$@H���    tH�D$@H�   H������H��8����������������H��HH�D$8����L��� A��   H��3 ��   ��\��H�D$ H�|$  tH�L$ �>���H�D$(�	H�D$(    H�D$(H�D$0H�D$0H��H�����������H�L$H��HH�D$PH�8 t>H�D$PH� H�D$(H�D$(H�D$ H�|$  t�   H�L$ �  H�D$0�	H�D$0    H�D$PH�     H��H��������������H�T$H�L$H��HH�D$PH�8 tH�� ��   ��  H�D$PH���    tH�� ��   ��  H�L$P�L���H�L$P�����H�D$PH�L$PH���   H�T$PH�°   H�T$0H�D$ L��H�D$PD���   H�T$XH�D$0H������H�L$P���   H�D$P���   uH�D$PH�8 uWH�D$PH�8 uH�D$P���   uH�D$Pǀ�   ����H�D$PH�     H�D$PH�   H������H�D$P���   ��   H�D$P���    ��   H�D$PH�   H�L$PH���   L��H��H�L$X��h ��u0H�D$Pǀ�       H�D$PW����   H��~ �  �  H�D$PH��H�T$XH��蜞��H�D$PH���D$     E3�A�   H��H�D$PH��2  H�L$P���   H�D$P���   tH�L$P����H�D$P���   �H�D$Pǀ�   ����H�D$P���   H��H��������������������H�L$H��(H�L$0�]���H�L$0�����H��(���������������L�D$�T$H�L$H��8H�D$@���    uH�D$@H���   ��   H�D$@���   9D$HuH�D$@H���   �   H�D$@H���L$H�L$ H�L$@L���   A�   H��H�D$@H��  H�L$@���   H�D$@���   u0H�D$@�L$H���   H�|$P tH�D$P�    H�D$@H���   �+H�D$@ǀ�   ����H�|$P tH�D$PH�L$@���   �3�H��8������������������H�T$H�L$H�|$ tH�D$H�L$���   � H�D$���    tH�D$���   �H�D$���   u�   �3�����������������������D�L$ L�D$H�T$H�L$H��HH��* H�@8H��$�   H�L$8��$�   �L$0H�L$xH�L$(�L$p�L$ D�L$hL�D$`H�T$XH�L$P�P(H��H��������H�T$H�L$H��(H�S* H�@8H�T$8H�L$0�PH��(����������������������H�L$H��(H�* H�@8H�L$0�PH��(����������������L�D$�T$H�L$H��(H��) H�@8L�D$@�T$8H�L$0�P H��(��������������H��(H��) H�@8�H��(�����������H�L$H��(H��) H�@8H�L$0H�	�PH�D$0H�     H��(�����������������D�L$ L�D$H�T$H�L$H��8H�L$@螏��H�D$ H�L$@菏��D�L$XL�D$PH�T$HH�H@H�D$ ���   H��8�������������D�L$ L�D$H�T$H�L$H��8H�L$@�>���H�D$ H�L$@�/���D�L$XL�D$PH�T$HH�H@H�D$ ���   H��8�������������H�L$H��8H�L$@����H���    u3��(H�L$@�Վ��H�D$ H�L$@�Ǝ��H�H@H�D$ ���   H��8�������������������L�L$ L�D$H�T$H�L$H��8H�L$@�~���H���    u3��7H�L$@�f���H�D$ H�L$@�W���L�L$XL�D$PH�T$HH�H@H�D$ ���   H��8���������������������L�L$ D�D$H�T$H�L$H��HH�L$P�����H���    u������?H�L$P����H�D$0H�L$P�ԍ���L$p�L$ L�L$hD�D$`H�T$XH�H@H�D$0���   H��H����������L�D$H�T$H�L$H��8H�L$@胍��H���    u������2H�L$@�h���H�D$ H�L$@�Y���L�D$PH�T$HH�H@H�D$ ���   H��8������������H�T$H�L$H��8H�L$@����H���    u������-H�L$@�����H�D$ H�L$@����H�T$HH�H@H�D$ ���   H��8����������������������L�D$H�T$H�L$H��   H�D$@����H��$�    tRH�L$H��S �H��$�   �~���H�D$8H��$�   �l���H�T$HH�H@H�D$8���   H��$�   �H�L$H�DT H��$�    tiH�L$`�R��H�D$0H�D$0H�D$(H�T$(H��$�   �^����H�L$`�S��H��$�   �����H���   H�D$ H�|$  tH�T$ H��$�   � ���H�Ĉ   ���������H�T$H�L$H��8H�L$@訋��H�D$ H�L$@虋��H�T$HH�H@H�D$ ���   H��8����������������̉T$H�L$H��8H�L$@�Y���H���    u� }  �,H�L$@�>���H�D$ H�L$@�/����T$HH�H@H�D$ ���   H��8��������L�L$ L�D$H�T$H�L$H��H�   �L$p�  ��t
�D$0   ��D$0    �T$0H�L$P�V����D$4H�L$`�dQ��;D$4H�L$`�,Q��;D$4~������?H�L$P葊��H�D$8H�L$P肊���L$p�L$ L�L$hL�D$`H�T$XH�H@H�D$8���   H��H��������L�L$ L�D$H�T$H�L$H��XH�L$`�.���H���    u������ZH�L$`����H�D$@H�L$`������$�   �L$0��$�   �L$(H��$�   H�L$ L�L$xL�D$pH�T$hH�H@H�D$@���   H��X���������������L�D$H�T$H�L$H��8H�L$@蓉��H���    u������2H�L$@�x���H�D$ H�L$@�i���L�D$PH�T$HH�H@H�D$ ���   H��8������������H�T$H�L$H��8H�L$@�(���H���    u�-H�L$@����H�D$ H�L$@����H�T$HH�H@H�D$ ���   H��8����������̉L$H��XH�L$0�~  H�T$0�L$`�J ��tH�|$0 u3�� �D$D�D$ D�L$@D�D$<�T$8H�L$0����H��X������������H�L$H��8H�D$@H� H�D$ H�L$ ��o��H�D$@H�     H��8����������������H�L$H��8H�D$@H� H�D$ H�L$ �o��H�D$@H�     H��8����������������H�L$H�D$������H�L$H��8H�D$@H��蚋���D$     �
�D$ ���D$ �|$ }HcD$ H�L$@H�D�(    ��H�D$@H��8�H�T$H�L$H��(H�D$0�     H�D$0H�@    H�! H��  E3�H�T$8H�L$0�PH�D$0H��(���H�L$H�D$H�     H�D$�@    H�D$�@    H�D$�@    H�D$�@    H�D$�@    H�D$��������������L�D$H�T$H�L$H�D$H�L$H�H�D$H�L$H�HH�D$�H�L$H��(H�D$0H���
���H��(������H�L$H��(H�(  H��  H�L$0�H��(��������������H�T$H�L$H�D$ÉT$�L$�D$�L$#ȋ������������̉T$H�L$H��(H�L$0������D$8����t
H�L$0�M��H�D$0H��(�����������H�T$H�L$H��8�   H�L$@�   H�D$ H�T$HH�L$ �  H�D$(3���tH�D$@H�@H��H�L$@H�AH�D$(H��8������H�T$H�L$H��8�   H�L$@�  H�й   ����H�D$ H�|$  t!H�L$H�_���H�L$ H� H�H�D$ H�D$(�	H�D$(    H�D$(H��8������H�T$H�L$H��XH�D$`H�@HD$hH�D$0H�D$`H�@H�L$`H�	H��H�D$(H�D$`H�@H9D$0��   A�   H�T$hH�D$`H�H�8  H�D$8H�D$8H��H�D$@H�L$`�  L�L$ H�L$@L��H�L$`H�H����  H�D$(H�|$( tp�D$ ��u3H�D$`H�8 t(H�D$`L�@H�T$(H�D$`H���  H�D$`H�������H�D$`H�L$(H�H�D$`H�L$8H�HH�D$`H�@H�L$(H��H�D$(�H�D$`H�@H�D$0H�D$`H�L$0H�HH�D$(H��X������������H�T$H�L$H��XH�D$`H�@HD$hH�D$0H�D$`H�@H�L$`H�	H��H�D$(H�D$`H�@H9D$0��   A�   H�T$hH�D$`H�H��   H�D$8H�D$8H��H�D$@H�L$`�k  L�L$ H�L$@L��H�L$`H�H����  H�D$(H�|$( tp�D$ ��u3H�D$`H�8 t(H�D$`L�@H�T$(H�D$`H���  H�D$`H������H�D$`H�L$(H�H�D$`H�L$8H�HH�D$`H�@H�L$(H��H�D$(�H�D$`H�@H�D$0H�D$`H�L$0H�HH�D$(H��X������������L�D$H�T$H�L$H��H�D$(H�L$ H�H��Hk�H�H+�H��H�$H�$H�H�|$0H��H�D$H�|$ uH�<$ uH�D$H�L$0H+�H��H�$H�H��H�$H�$H�������H�T$H�L$H��8H�T$@�   ����H�D$ H�|$  tH�D$ H�L$HH�	H�H�D$ H�D$(�	H�D$(    H�D$(H��8��������H�L$H��H�D$ H�8 t&H�D$ H�@H��H�$�H�$H��H�$H�<$ |��H�D$ H�@    H�������H�L$H��H�D$ H�8 t&H�D$ H�@H��H�$�H�$H��H�$H�<$ |��H�D$ H�@    H�������H�L$H�D$H�@��H�L$H�D$������H�L$H�D$������H�L$H�D$H� ���H�L$H�D$H�@H%��� ������������H�L$H��(H�8 H��  H�L$0�PpH��(�������������L�D$H�T$H�L$H��(H�D$@H��L��H�T$0H�L$8�� H��(�������������L�D$H�T$H�L$H��(H�D$@H��L��H�T$0H�L$8��� H��(�������������L�D$H�T$H�L$H��8H�L$P����H�D$ H�L$P����H�e H�IH�L$(H�T$ L��D���T$HH�L$@H�D$(��0  H��8�L�L$ L�D$H�T$H�L$H��8H�D$X� A��   H�#l H�L$ �y���L��H�T$PH�L$H�W���H��8���L�L$ L�D$H�T$H�L$H��8H�D$X� A��   H��k H�L$ �)���L��H�T$PH�L$H����H��8���H�T$�L$H��(H�� H�@H�T$8�L$0��`  H��(�����H�L$H�D$H�s H�H�D$H�@    H�D$H�@    H�D$�@    H�D$�����������������H�L$H��(H�D$0H��r H�H�D$0�x uH�� H�@hH�L$0H�I�H�D$0H�@    H�D$0H�@    H��(���������H�L$�   ����������������������H�L$�   ����������������������L�D$H�T$H�L$3����������������D�D$�T$H�L$������������������D�L$ D�D$�T$H�L$H��8��  H�L$@�:  �D$`�D$ D�L$XD�D$P�T$HH�L$@�:  2�H��8��������������������D�L$ D�D$�T$H�L$H��8H�D$@H� �L$`�L$ D�L$XD�D$P�T$HH�L$@�P(H��8���������������H�T$H�L$3���������������������L�D$�T$H�L$�   �������������H�T$H�L$����������������������L�D$H�T$H�L$H��h�D$4    H�L$x�k�  �D$0�|$0INIbG�|$0INIbtv�|$0$'  ��  �|$0MicM��  �|$0SACb��   �|$0ARDb�  �  �|$0NPIb��  �|$0ISIb��   �|$0NIVbt0�|$0cnys��  ��  H�D$pH� H�L$p�P�D$4   �  H�D$pH� H�L$p�P�D$4   �  �D$<    �D$8    H�D$pH� L�D$8H�T$<H�L$p�P��t H� H�@hD�D$8�T$<H�L$pH�I�P(�D$4   �A  H�L$p��  �D$TH�L$p�  H�L$pH�	H�L$X�T$TD��H�L$pH�D$X�P �D$4   ��   E3��   H�L$x�;A���D$HE3��   H�L$x�%A���D$DE3��   H�L$x�A���D$LE3��   H�L$x��@���D$@H�D$pH� H�L$xH�L$(�L$@�L$ D�L$LD�D$D�T$HH�L$p�P0�D$4   �gH�D$pH� H�T$xH�L$p�P8�TH�D$pH� H�T$xH�L$p�PH�D$4   �1E3��IicMH�L$x�s@���D$PH�D$pH� L�D$x�T$PH�L$p�P@��D$4H��h��������������̉T$H�L$H��   H�D$@����H��$�   H�x ��   ��$�    tFH��$�   ��   �D$ H��$�   H�I����H�) H�I`H�L$8�T$ H��H�D$8���   �lH��$�   �   ��H�L$X�+�  �ARDbH�L$h��@ H�D$0H�D$0H�D$(L�L$(L�D$XH�T$HH��$�   H�H�}  H�L$H�s����H�L$h�A H�Ĉ   �����������������H�T$H�L$H��(H�s H�@hH�T$8H�L$0H�I���   �   H��(����������H�L$H��(H�8 H�@hH�L$0H�I�P H��(������������H�L$H��(H� H�@hH�L$0H�I�PH��(������������H�L$H��(H�� H�@hH�L$0H�I�PH��(������������H�L$H��(H�� H�@hH�L$0H�I���   H��(���������H�L$H��(H�x H�@hH�L$0H�I���  H��(��������̉T$H�L$H��(H�D H�@h�T$8H�L$0H�I�PPH��(��������������������L�L$ D�D$�T$H�L$H��(H�� H�@hL�L$HD�D$@�T$8H�L$0H�I�PXH��(����������������L�D$�T$H�L$H��(H�� H�@hL�D$@�T$8H�L$0H�I�P`H��(����������H�L$H��(H�x H�@hH�L$0H�I�PhH��(�����������̉T$H�L$H��(H�D H�@h�T$8H�L$0H�I���  H��(�����������������H�T$H�L$H��(H� H�@hH�T$8H�L$0H�I�P@H��(�����������������̉T$H�L$H��(H�� H�@h�T$8H�L$0H�I�PHH��(��������������������H�T$H�L$H��(H�L$8��  ��uH�L$8�i�  H��H�L$0�L����8H�L$8���  ��uH�L$8������H�L$0�e����H�,c �
  ����H��(��������������D�D$�T$H�L$H��(H�� H�@hD�D$@�T$8H�L$0H�I���   H��(�������D�D$H�T$H�L$H��(H�� H�@hD�D$@H�T$8H�L$0H�I���   H��(���������������������L�D$�T$H�L$H��(H�o H�@hL�D$@�T$8H�L$0H�I���   H��(�������L�D$H�T$H�L$H��(H�. H�@hL�D$@H�T$8H�L$0H�I���   H��(���������������������L�D$H�T$H�L$H��hH�L$x�C�  ����   H��$�   �-�  ��uMH��$�   諛  H�D$(H�L$x蜛  H�� H�IhH�L$0H�T$(L��H��H�D$pH�HH�D$0���   �nH��$�   �Κ  ��uKH��$�   �����D$ H�L$x�>�  H�? H�IhH�L$8�T$ D��H��H�D$pH�HH�D$8���   �H�'a ��  �m�����   H�L$x�^�  ����   H��$�   �H�  ��uLH��$�   �ƚ  H�D$@H�L$x�w���H�� H�IhH�L$HH�T$@L��H�D$pH�HH�D$H���   �mH��$�   ��  ��uJH��$�   �(����D$$H�L$x����H�[ H�IhH�L$P�T$$D��H�D$pH�HH�D$P���   �H�d` ��  �����H�q` ��  �w���H��h�������������������L�L$ L�D$�T$H�L$H��8H�� H�@`H�L$`H�L$ L�L$XL�D$P�T$HH�L$@H�I���  H��8������������������̉T$H�L$H��(H�� H�@`�T$8H�L$0H�I���  H��(������������������\$ D�D$�T$H�L$H��(H�9 H�@`�\$HD�D$@�T$8H�L$0H�I���  H��(�����������D�L$ D�D$�T$H�L$H��8H��
 H�@h�L$`�L$ D�L$XD�D$P�T$HH�L$@H�I�P0H��8��������D�L$ D�D$�T$H�L$H��8H��
 H�@h�L$`�L$ D�L$XD�D$P�T$HH�L$@H�I�P8H��8��������D�L$ D�D$H�T$H�L$H��hH�I
 H�@h��$�   �L$P��$�   �L$H��$�   �L$@��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ D��$�   D��$�   H�T$xH�L$pH�I���   H��h��������D�L$ D�D$H�T$H�L$H��8H��	 H�@h�L$`�L$ D�L$XD�D$PH�T$HH�L$@H�I��  H��8�������������������L�L$ �T$�L$H�L$H��HH�G	 H�@h��$�   �L$0�L$x�L$(�L$p�L$ L�L$h�T$`�L$XH�L$PH�I��0  H��H������������D�L$ D�D$H�T$H�L$H��h�D$P�����D$H�����D$@������$�   �D$8��$�   �D$0�D$(�����D$ ����A�����A�����H�T$xH�L$p����H��h����������̉T$H�L$H��(H�d H�@h�T$8H�L$0H�I�PpH��(��������������������H�T$H�L$H��(H�# H�@hH�T$8H�L$0H�I�PxH��(������������������D�D$H�T$H�L$H��(H�� H�@hD�D$@H�T$8H�L$0H�I���  H��(���������������������H�L$H��(H�� H�@hH�L$0H�I���   H��(���������H�L$H��(H�h H�@hH�L$0H�I��  H��(����������L$H�L$H��(H�2 H�@h�L$8H�L$0H�I��  H��(�������������D�L$ D�D$�T$H�L$H��8H�� H�@h�L$`�L$ D�L$XD�D$P�T$HH�L$@H�I���   H��8���������������������H�L$H��(H�� H�@hH�L$0H�I���   H��(���������H�L$H��(H�h H�@hH�L$0H�I���   H��(���������D�L$ D�D$�T$H�L$H��8H�* H�@h�L$`�L$ D�L$XD�D$P�T$HH�L$@H�I��   H��8���������������������D�L$ D�D$�T$H�L$H��HH�� H�@h��$�   �L$0�L$x�L$(�L$p�L$ D�L$hD�D$`�T$XH�L$PH�I���   H��H������������������L�D$H�T$H�L$H��(H�^ H�@hL�D$@H�T$8H�L$0H�I��   H��(���������������������L�D$H�T$H�L$H��(H� H�@hL�D$@H�T$8H�L$0H�I���   H��(���������������������L�D$H�T$H�L$H��(H�� H�@hL�D$@H�T$8H�L$0H�I��(  H��(���������������������L�D$H�T$H�L$H��(H�n H�@hL�D$@H�T$8H�L$0H�I���   H��(���������������������H�L$H��XH�D$0�����YALfH�L$8��1 H�D$ H�D$ H�D$(H�T$(H�L$`�q����H�L$8�V2 H��X������������������L�L$ L�D$H�T$H�L$H��(H�|$@ tE3��   H�L$8�[0��H�L$@�H�|$H tE3��   H�L$8�:0��H�L$H�H�w H�@hL�D$HH�T$@H�L$0H�I���   H��(��������������L�L$ L�D$H�T$H�L$H��(L�L$HL�D$@H�T$8H�D$0H�H�+K  H��(�������L�L$ D�D$H�T$H�L$H��8H�� H�@h�L$`�L$ L�L$XD�D$PH�T$HH�L$@H�I���   H��8������������������̉T$H�L$H��(H�� H�@h�T$8H�L$0H�I���   H��(�����������������L�L$ L�D$�T$H�L$H��8H�J H�@hH�L$hH�L$(H�L$`H�L$ L�L$XL�D$P�T$HH�L$@H�I��   H��8���������D�L$ D�D$�T$H�L$H��8H�� H�@h�L$h�L$(�L$`�L$ D�L$XD�D$P�T$HH�L$@H�I��  H��8�������������D�L$ D�D$H�T$H�L$H��x�D$0    �D$4    L�L$8L�D$<H��$�   H��$�   H�H��H  H��$�   ������H�L$X�|�  H�D$HH�D$(H�D$DH�D$ L�L$4L�D$0H�T$XH��$�   H�H�H  ��$�    t\��$�    tR�D$09D$<~8�D$D�L$0ȋ�9D$<}&�D$49D$8~�D$H�L$4ȋ�9D$8}
�D$@   ��D$@    �D$@�r�>��$�    t4�D$49D$8~�D$H�L$4ȋ�9D$8}
�D$P   ��D$P    �D$P�2�D$09D$<~�D$D�L$0ȋ�9D$<}
�D$L   ��D$L    �D$LH��x���������������\$ �T$�T$H�L$H��8H�  H�@h�L$`�L$ �\$X�T$P�T$HH�L$@H�I���  H��8�����������������L�L$ L�D$H�T$H�L$H��(H��� H�@hL�L$HL�D$@H�T$8H�L$0H�I���  H��(�����������H�L$H��(H�h� H�@hH�L$0H�I���  H��(���������H�L$H��(H�8� H�@hH�L$0H�I��8  H��(���������H�L$H��(H�D$0H�#Z H�H��� H�@`H�T$0H��u  �H�L$0H�AH�D$0�@    H�D$0H��(�����������������H�L$H��(H�D$0H��Y H�H�D$0H�x tH��� H�@`H�L$0H�I�PH�D$0H�@    H��(��������������������H�L$�   ����������������������H�L$�   ����������������������L�D$�T$H�L$�   �������������L�D$�T$H�L$3�����������������H�L$3����������H�T$H�L$����������������������H�L$�����������L�D$H�T$H�L$H��8H�L$H��  �D$ �|$ NIVbG�|$ NIVb��   �|$ $'  ��  �|$ MicM�  �|$ TCAb�4  �|$ INIbtD�  �|$ ckhc�P  �|$ ytsdt]�|$ atnit�|$ cnys��   �Y  �; �O  H�D$@�x t
�   �<  H�D$@�@   H�D$@H� H�L$@�P�  H�D$@H� H�L$@�P8H�D$@�@    ��   H�D$@�x u
�   ��   H�D$@H� H�L$@�P��   E3��IicMH�L$H�	)���D$$H�D$@H� L�D$H�T$$H�L$@�P�   E3��IicMH�L$H��(���D$$H�D$@H� L�D$H�T$$H�L$@�P�kE3��diemH�L$H�(���D$$H�D$@H� L�D$H�T$$H�L$@�P �D$(�D$(�2H�D$@H� H�L$@�P(� �H�D$@H� H�T$HH�L$@�P0�   �3�H��8����������D�L$ D�D$�T$H�L$H��XH�D$`H�x u3��   H�W� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    ��$�   �L$ E3�D�D$p�   H�L$`H�I��  H��� H�@`��$�   �L$0��$�   �L$(��$�   �L$ D�L$xE3��T$hH�L$`H�I��0  H��X���������������H�L$H��(H�D$0H�x u3��H��� H�@`H�L$0H�I�PH��(�����������̉T$H�L$H��(H�L$0����H��(���������������������L�L$ L�D$H�T$H�L$H��xH�D$X�����D$0    H��$�   H�x u(3�H��$�   �Y{  ��D$0���D$0H��$�   �   H��$�   �s�  H�D$8H��$�   �!�  H��� H�I`H�L$@H�T$8H�T$ L��$�   D��H��$�   H�PH�L$`H�D$@���  H�D$HH�D$HH�D$PH�T$PH��$�   �����D$0���D$0H�L$`�
���H��$�   H��x��������������H�T$H�L$H��(H�� H�@`H�T$8H�L$0H�I��(  H��(���������������H�L$H��8H�L$@�-���H��� H�I`H�L$ H��H�D$ ��  H��8�����������H�L$H��XH��� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��4   H�L$`H�I��  H��X������������H�L$H��XH�(� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��;   H�L$`H�I��  H��X�����������̉T$H�L$H��(H��� H�@`�T$8H�L$0H�I�P(H��(��������������������H�T$H�L$H��XH�D$`H�x u�YH�e� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     L�L$hE3��   H�L$`H�I��  H��X�������L�L$ D�D$�T$H�L$H��(H��� H�@hL�L$HD�D$@�T$8H�L$0H�I�PXH��(����������������L�D$�T$H�L$H��(H��� H�@hL�D$@�T$8H�L$0H�I�P`H��(����������H�L$H��(H�h� H�@hH�L$0H�I�PhH��(������������D�D$H�T$H�L$H��8H�D$@H�x u3��IH�L$H�Ä  H�D$ H�L$H�t�  H�� H�I`H�L$(H�T$ L��D�D$P��H�D$@H�HH�D$(�P H��8����������������H�T$H�L$H��8H�D$@H�x u3��GH�L$H�H�  H�D$ H�L$H���  H��� H�I`H�L$(H�T$ L��H�D$@H�HH�D$(���  H��8�������D�L$ D�D$H�T$H�L$H��h��$�    u
�D$P   ��D$P   �D$@����D$8  ���$�   �D$0�D$(    �D$P�D$ E3�D��$�   H�T$xH�L$p�   H��h�������������������D�L$ D�D$H�T$H�L$H��xH�D$8�����tnivH�L$P�" �D��$�   �ulavH�L$P�S!��A�gnlf�tmrfH�L$P�>!��D��$�   �inimH�L$P�'!��D��$�   �ixamH�L$P�!��D��$�   �petsH�L$P�� ��D��$�   �sirtH�L$P�� ����$�     �u��$�   ���t.D��$�   �2nimH�L$P� ��D��$�   �2xamH�L$P� ��L�L$PL��$�   H�T$@H��$�   �p���H�D$(H�D$(H�D$0H�L$0�G����D$ H�L$@�I����H�L$P��! �D$ H��x�����������������������\$ �T$H�T$H�L$H��xH�D$8�����tlfvH�L$P�! ���$�   �ulavH�L$P�Ղ  D��$�   �tmrfH�L$P������$�   �inimH�L$P覂  ��$�   �ixamH�L$P莂  ��$�   �petsH�L$P�v�  D��$�   �sirtH�L$P�j����$�   f.>O zu��$�   f.)O zt0��$�   �2nimH�L$P��  ��$�   �2xamH�L$P��  D��$�   �dauqH�L$P����L�L$PL��$�   H�T$@H��$�   �����H�D$(H�D$(H�D$0H�L$0�����D$ H�L$@�����H�L$P�=  �D$ H��x����������������������\$ �T$H�T$H�L$H��h��$�   �D$P�D$H    W��D$@W��D$8�D$0temf��$�   �D$(��$�   �D$ ��$�   ��$�   H�T$xH�L$p�����H��h�����������������������\$ �T$H�T$H�L$H��x��$�   f.�M zu��$�   �D$`���$�   �  �D$`��$�   f.�M zu��$�   �D$h���$�   �H  �D$h��$�   �4  ��$�   �D$P�D$H    W��L$@W��L$8�D$0rgdf�D$(�D$`�D$ �\$h��$�   H��$�   H��$�   �����H��x��������������\$ �T$H�T$H�L$H��h��$�   �^�L ��$�   �^�L ��$�   �^�L ��$�   �D$P�D$H    W��\$@W��\$8�D$0tcpf�D$(�L$ (���$�   H�T$xH�L$p����H��h�����������L�L$ L�D$H�T$H�L$H��   H�D$h����H��$�    uH�"� H�@��0  H��$�   H��$�    u3���  H��$�   ��o �D$ �tlfvH�L$(�� �H��$�   �z  �*L$ �Y��)x  �D$PH��$�   �fy  �x  �L$P�^�(�(кulavH�L$(�R~  A�mrff�tmrfH�L$(�H��H��$�   �0z  �*L$ �Y���w  �D$XH��$�   ��x  �w  �L$X�^�(�(кinimH�L$(��}  H��$�   ��y  �*L$ �Y��nw  �D$@H��$�   �x  �Vw  �L$@�^�(�(кixamH�L$(�}  ��7 �petsH�L$(�}  E3��dauqH�L$(�y��D�D$ �spffH�L$(�e��D��$�   �sirtH�L$(�N��L�L$(L��$�   H�T$pH��$�   �$���H�D$`H�D$`H�D$HH�L$H������D$$H�L$p������H�L$(� �D$$H�Ĉ   �������D�L$ L�D$H�T$H�L$H��xH�D$8�����CITbH�L$P�� �L��$�   �CITbH�L$P�%��D��$�   �sirtH�L$P���D��$�   �ulavH�L$P�u��L�L$PL��$�   H�T$@H��$�   �K���H�D$(H�D$(H�D$0H�L$0�"����D$ H�L$@�$����H�L$P� �D$ H��x������������������\$ L�D$H�T$H�L$H��XH�D$`H�x u3��kH�L$h�z  H�D$@H�L$h�^z  H��� H�I`H�L$HH�T$@H�T$0��$�   �T$(��$�   �D$ �\$xL�D$p��H�D$`H�HH�D$H�PPH��X��������D�L$ L�D$H�T$H�L$H��xH�D$H����H�T$PH��$�   �=X��H�D$8H�D$8H�D$@�D$     D��$�   L�D$@H��$�   H��$�   �����D$0H�L$P����D$0H��x��������������L�D$H�T$H�L$H��HH�D$PH�x u3��uH�L$X�y  H�D$0H�L$X�4y  H��� H�I`H�L$8H�T$0L��L�D$$��H�D$PH�HH�D$8�PX�D$(�|$$ t
�D$    ��D$     H�D$`�L$ ��D$(H��H��������������������L�D$H�T$H�L$H��8H�D$@H�x u3��IH�L$H��x  H�D$ H�L$H�x  H�� H�I`H�L$(H�T$ L��L�D$P��H�D$@H�HH�D$(�PXH��8����������������L�D$H�T$H�L$H��8H�D$@H�x u3��IH�L$H�Sx  H�D$ H�L$H�x  H��� H�I`H�L$(H�T$ L��L�D$P��H�D$@H�HH�D$(�P`H��8����������������L�L$ L�D$H�T$H�L$H��(H�D$PL��H�T$8H�L$0�Q�����u3��KH�D$PH��L��H�T$@H�L$0�.�����u3��(H�D$PH��L��H�T$HH�L$0������u3���   H��(����������L�D$H�T$H�L$H��hH�D$pH�x u3���   H�D$(    H�L$x�7w  H�D$8H�L$x��v  H�y� H�I`H�L$@H�T$8L��L�D$(��H�D$pH�HH�D$@�Pp�D$ �|$  tfH�|$( t^H�T$(H��$�   ����H�|$( t;H�D$(H�D$HH�D$HH�D$0H�|$0 t�   H�L$0�m  H�D$P�	H�D$P    H�D$(    �D$ H��h���������������L�L$ L�D$H�T$H�L$H��HH�D$PH�x u3��PH�L$X�>v  H�D$0H�L$X��u  H��� H�I`H�L$8H�T$0H�T$ L�L$hL�D$`��H�D$PH�HH�D$8�PxH��H��������������������L�L$ L�D$H�T$H�L$VWH��HH�|$p uH�� H�@��0  H�D$pH�|$p u3��bH�L$p��g �D$ L�D$(H�T$hH�L$`������D$$�*D$ �Y�C �L$(�Y�C (�H�L$0�L H�|$xH��   �D$$H��H_^��������������������L�D$H�T$H�L$H��XH�D$0����H�L$8�H���L�D$8H�T$hH�L$`�u����D$ �|$  u�D$$    H�L$8����D$$�%H�T$8H�L$p�cS���D$ �D$(H�L$8�l���D$(H��X���������H�T$H�L$H��hH�D$pH�x u3��{H�L$x�ht  H�D$PH�L$x�t  H��� H�I`H�L$XH�T$PH�T$HH�D$@    �D$8    �D$0    �D$(    �D$     E3�D���1   H�D$pH�HH�D$X��  H��h�������������������D�L$ L�D$H�T$H�L$H��(E3��T$HH�L$@�n  E3�D��H�T$8H�L$0����H��(��������������D�L$ L�D$H�T$H�L$H��XE3��T$xH�L$p�t����$�   �L$@��$�   �L$8�D$0    ��$�   �L$(��$�   �L$ D��$�   D��H�T$hH�L$`����H��X���������������������D�L$ L�D$H�T$H�L$H��hWҋ�$�   H��$�   �p  �D$P    ��$�   �D$H��$�   �L$@��$�   �L$8��$�   �D$0��$�   �L$(��$�   �L$ ��$�   (�H�T$xH�L$p�\���H��h��������D�L$ L�D$H�T$H�L$H��HWҋT$hH�L$`�Wo  �D$0    ��$�   �L$(�L$x�L$ �\$p(�H�T$XH�L$P����H��H��������D�L$ L�D$H�T$H�L$H��HWҋT$hH�L$`��n  �D$0    ��$�   �L$(�L$x�L$ �\$p(�H�T$XH�L$P����H��H��������D�L$ L�D$H�T$H�L$H��HWҋT$hH�L$`�wn  �D$0    ��$�   �L$(�L$x�L$ �\$p(�H�T$XH�L$P�\���H��H��������L�L$ L�D$H�T$H�L$H��hH�L$@�>c  L��D��$�   H�T$PH��$�   �1n  �D$8    ��$�   �L$0H��$�   H�L$(H��$�   H�L$ L��L��$�   H�T$xH�L$p�z���H��h����������������������D�L$ L�D$H�T$H�L$H��   H�D$X����H�L$x���H�D$HH�D$HH�D$PL�L$PD��$�   H�T$`H��$�   ��E��H�D$8H�D$8H�D$@��$�   �D$ E3�L�D$@H��$�   H��$�   �����D$0H�L$`����H�L$x����D$0H�Ę   ���������D�L$ L�D$H�T$H�L$H��   H�D$H����H�L$x��J��H�D$8H�D$8H�D$@L�L$@D��$�   H�T$PH��$�   �dk  H�D$(H�D$(H�D$0E3�L�D$0H��$�   H��$�   ������D$ H�L$P�*L���H�L$x�L���D$ H�Ĩ   ��������������������D�L$ L�D$H�T$H�L$H��x�* �D$0��$�   �tWҋ�$�   H��$�   ��k  �D$0H�L$8�1��L��D��$�   H�T$PH��$�   �����$�   �L$(��$�   �D$ �\$0L��H��$�   H��$�   �T���H��x����������������D�L$ L�D$H�T$H�L$H��8�D$     L�D$ H�T$HH�L$@�<����D$$D�D$ �T$XH�L$P�n  �D$$H��8�������������D�L$ L�D$H�T$H�L$H��8L�D$ H�T$HH�L$@�����D$$D�D$ �T$XH�L$P����D$$H��8���������������������D�L$ L�D$H�T$H�L$H��8L�D$(H�T$HH�L$@�����D$ �T$(�T$XH�L$P�<n  �D$ H��8��������������������L�L$ L�D$H�T$H�L$H��HH�L$(�>_  L�L$(L�D$`H�T$XH�L$P������D$ L�D$(�T$pH�L$h�n  �D$ H��H����������������������L�L$ L�D$H�T$H�L$H��HH�L$ ���L�D$ H�T$XH�L$P�������u3��PL�D$(H�T$`H�L$P������u3��4L�D$0H�T$hH�L$P������u3��L�D$ �T$xH�L$p� 
���   H��H��������������D�L$ L�D$H�T$H�L$H��XH�D$(����H�L$0�
���L�D$0H�T$hH�L$`�@����D$ L�D$0�T$xH�L$p�F
���D$ �D$$H�L$0�R
���D$$H��X���������������D�L$ L�D$H�T$H�L$H��hH�D$(����H�L$0��F���L�D$0H�T$xH�L$p�����D$ L�D$0��$�   H��$�   ��k  �D$ �D$$H�L$0�!H���D$$H��h���������D�L$ L�D$H�T$H�L$H��XH�L$0�v	��L�L$(L�D$0H�T$hH�L$`�E����D$ �|$x�tL�D$0�T$xH�L$p�����$�   �t�T$(��$�   H�L$p�k  �D$ H��X��������������L�D$H�T$H�L$H��8H�L$P�3i  � �D$$H�L$P�h  �D$ �|$  t�D$$   D�L$ D�D$$H�T$HH�L$@����H��8�������������������D�L$ L�D$H�T$H�L$H��hH��$�   ��g  �D$PH��$�   �h  ��$�   �L$@��$�   �L$8�L$P�L$0��$�   �L$(��$�   �L$ D��$�   D� H�T$xH�L$p�����H��h���������\$ L�D$H�T$H�L$H��xH��$�   �jg  �D$`H��$�   �9h  �L$`�L$P��$�   �L$H��$�   �D$@��$�   �D$8��$�   �L$0��$�   �D$(��$�   �D$ ��$�   �H��$�   H��$�   ����H��x����������\$ L�D$H�T$H�L$H��XH�L$p�f  �D$@H�L$p�g  �L$@�L$0��$�   �D$(��$�   �D$ �\$x�H�T$hH�L$`�����H��X�������������\$ L�D$H�T$H�L$H��XH�L$p�-f  �D$@H�L$p��f  �L$@�L$0��$�   �D$(��$�   �D$ �\$x�H�T$hH�L$`�����H��X�������������\$ L�D$H�T$H�L$H��XH�L$p�e  �D$@H�L$p�f  �L$@�L$0��$�   �D$(��$�   �D$ �\$x�H�T$hH�L$`����H��X������������L�L$ L�D$H�T$H�L$H��XH�L$x�^e  �D$@H�L$x� f  �L$@�L$8��$�   �L$0H��$�   H�L$(H��$�   H�L$ L��L�D$pH�T$hH�L$`����H��X��������D�L$ L�D$H�T$H�L$H��HH�L$`�e  �D$0H�L$`�e  �L$h�L$ �L$0D��L��H�T$XH�L$P����H��H�����������D�L$ D�D$H�T$H�L$H��   H�D$p�����gnrsH�L$8�M ���$�   H�L$P��X  �L�D$P�   H�L$8�Vf  �H�L$P�������$�   H�L$`�X  �L�D$`�   H�L$8�%f  �H�L$`�ʶ��L�L$8L��$�   H�T$xH��$�   ����H�D$0H�D$0H�D$(H�L$(肼���D$ H�L$x脶���H�L$8� �D$ H�Ę   ���������������\$ L�D$H�T$H�L$H��8H�L$P�=d  �L$h�L$(�D$`�D$ �\$XL��H�T$HH�L$@����H��8�������������H�L$H��XH�(� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��    H�L$`H�I��  H��X������������L�D$H�T$H�L$H��(H�D$0H�x u3��$H��� H�@hL�D$@H�T$8H�L$0H�I��   H��(���������������������L�D$H�T$H�L$H��(H�D$0H�x u3��$H�>� H�@hL�D$@H�T$8H�L$0H�I���   H��(���������������������L�D$H�T$H�L$H��(H�D$0H�x u3��$H��� H�@hL�D$@H�T$8H�L$0H�I���   H��(���������������������L�D$H�T$H�L$H��(H�D$0H�x u3��$H�~� H�@hL�D$@H�T$8H�L$0H�I��(  H��(���������������������L�L$ L�D$�T$H�L$H��HH�L$P����H� � H�I`H�L$0H�T$pH�T$ L�L$hL�D$`�T$XH��H�D$0���  H��H���������������������D�L$ D�D$H�T$H�L$H��hH�L$x�^b  H�D$PH�L$x�b  H��� H�I`H�L$XH�T$PH�T$HH�D$@    �D$8    �D$0    ��$�   �T$(��$�   �T$ E3�D���=   H�D$pH�HH�D$X��  H��h�������������������L�L$ D�D$H�T$H�L$H��hH�L$x�a  H�D$PH�L$x�_a  H��� H�I`H�L$XH�T$PH�T$HH��$�   H�T$@�D$8    �D$0    �D$(������$�   �T$ E3�D���=   H�D$pH�HH�D$X��  H��h������������������D�L$ L�D$�T$H�L$H��8H�|$P uH�� H�D$PH�L$P�6��H�<� H�I`H�L$ D�L$XL���T$HH�D$@H�HH�D$ ���   H��8�������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��vH�D$P    H��� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ L��$�   D�D$x�   H�L$pH�I��  H�D$PH��h���������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��vH�D$P    H�!� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ L��$�   D�D$x�   H�L$pH�I��  H�D$PH��h���������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��yH�D$P    H�q� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ L��$�   D�D$x�   H�L$pH�I��  H�D$PH��h������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��tH�D$P    H��� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h�����������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��tH�D$P    H�� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h�����������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��tH�D$P    H�a� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�*   H�L$pH�I��  H�D$PH��h�����������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��qH�D$P    H��� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h��������������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��qH�D$P    H�� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h��������������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��qH�D$P    H�Q� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�	   H�L$pH�I��  H�D$PH��h��������������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��qH�D$P    H��� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�
   H�L$pH�I��  H�D$PH��h��������������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��tH�D$P    H��� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h�����������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��tH�D$P    H�A� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h�����������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��vH�D$P    H��� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ L��$�   D�D$x�'   H�L$pH�I��  H�D$PH��h���������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��vH�D$P    H��� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ L��$�   D�D$x�,   H�L$pH�I��  H�D$PH��h���������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��tH�D$P    H�1� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�:   H�L$pH�I��  H�D$PH��h�����������������D�D$�T$H�L$H��hH�D$pH�x u3��iH�D$P    H��� H�@`H�L$PH�L$HH�D$@    �D$8    �D$0    �L$x�L$(��$�   �L$ E3�E3��)   H�L$pH�I��  H�D$PH��h�����������������D�D$�T$H�L$H��hH�D$pH�x u3��iH�D$P    H��� H�@`H�L$PH�L$HH�D$@    �D$8    �L$x�L$0�D$(    ��$�   �L$ E3�E3��)   H�L$pH�I��  H�D$PH��h�����������������D�L$ D�D$�T$H�L$H��XH�D$`H�x u3��\H�J� H�@`H�D$H    H�D$@    �D$8    ��$�   �L$0�L$x�L$(�L$p�L$ E3�D�D$h�   H�L$`H�I��  H��X���������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��tH�D$P    H��� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h�����������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��tH�D$P    H�� H�@`H�L$PH�L$HH�D$@    ��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�>   H�L$pH�I��  H�D$PH��h�����������������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��qH�D$P    H�Q� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h��������������������D�L$ D�D$�T$H�L$H��XH��� H�@`H�D$H    H�D$@    �D$8    ��$�   �L$0�L$x�L$(�L$p�L$ E3�D�D$h�.   H�L$`H�I��  H��X���������L�L$ D�D$H�T$H�L$H��hH�D$pH�x u3��   H�L$x��Q  H�D$PH�L$x�|Q  H�� H�I`H�L$XH�T$PH�T$HH�D$@    �D$8    �D$0    �D$(    ��$�   �T$ L��$�   D���   H�D$pH�HH�D$X��  H��h��������������H�T$H�L$H��hH�D$pH�x u3��{H�L$x�Q  H�D$PH�L$x��P  H�Z� H�I`H�L$XH�T$PH�T$HH�D$@    �D$8    �D$0    �D$(    �D$     E3�D���   H�D$pH�HH�D$X��  H��h�������������������L�D$H�T$H�L$H��8H�D$@H�x u3��LH�L$H�cP  H�D$ H�L$H�P  H��� H�I`H�L$(H�T$ L��L�D$P��H�D$@H�HH�D$(���   H��8�������������L�D$H�T$H�L$H��HH�T$`H�L$0�.�  L�D$(H�T$ H�L$0��  ��t5H�|$( u��H�L$(�R&��L��D�D$ H�T$XH�L$P������u3��본   H��H��������D�L$ D�D$�T$H�L$H��hH�D$pH�x u3��qH�D$P    H��� H�@`H�L$PH�L$HH�D$@    �D$8    ��$�   �L$0��$�   �L$(��$�   �L$ E3�D�D$x�   H�L$pH�I��  H�D$PH��h��������������������D�L$ L�D$H�T$H�L$H��XH�� H�@hH�L$hH�I�H�D$hH�@    H�D$hH�L$`H�HH�L$p�N  H�D$8H�L$p�>N  H�Ͽ H�I`H�L$@H�T$8H�T$ D�L$xL�D$h��H�D$`H�HH�D$@��8  H�L$hH�AH�D$hH�x t
�D$0   ��D$0    �D$0H��X���������������������D�L$ D�D$�T$H�L$H��XH�D$`H�x u3��\H�*� H�@`H�D$H    H�D$@    �D$8    ��$�   �L$0�L$x�L$(�L$p�L$ E3�D�D$h�/   H�L$`H�I��  H��X���������D�D$H�T$H�L$H��8H�|$H u3��OH�D$H�@    H�L$H����H�D$ H�L$@�ܣ��H�}� H�I`H�L$(H�T$ L�T$PH��H�D$(��   H��8�������������̉T$H�L$H��XH�D$`H�x u3��WH�$� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �L$h�L$ E3�E3��   H�L$`H�I��  H��X��������H�L$H��hH�L$p����H��� H�I`H�L$PH�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��6   H��H�D$P��  H��h��������������D�L$ D�D$�T$H�L$H��(H�D$0H�x u3��(H�� H�@`D�L$HD�D$@�T$8H�L$0H�I���   H��(�������������D�L$ D�D$�T$H�L$H��XH�D$`H�x u3��aH��� H�@`��$�   �L$@��$�   �L$8��$�   �L$0H��$�   H�L$(��$�   �L$ D�L$xD�D$p�T$hH�L$`H�I���  H��X��������������������H�L$H��(H�D$0H�x u3��H�(� H�@`H�L$0H�I���   H��(���������D�D$�T$H�L$H��(H�D$0H�x u3��#H�߻ H�@`D�D$@�T$8H�L$0H�I���   H��(������̉T$H�L$H��8H�D$@H�x u3��.�D$H��H��� H�I`H�L$ ��H�D$@H�HH�D$ ���   H��8����������������̉T$H�L$H��(H�D$0H�x u3��H�4� H�@`�T$8H�L$0H�I���   H��(�����������������D�L$ D�D$�T$H�L$H��8H�D$@H�x u3��0H�ں H�@`�L$`�L$ D�L$XD�D$P�T$HH�L$@H�I���   H��8���������������������L�D$H�T$H�L$H��   H�D$h����H�L$p��  �H��$�   �	I  H�D$XH��$�   �H  H�H� H�I`H�L$`H�T$XH�T$HH�T$pH�T$@�D$8    �D$0    �D$(    �D$     E3�D���8   H��$�   H�HH�D$`��  �D$P�|$P tH�T$pH��$�   �T�  �D$P�D$TH�L$p�"�  �D$TH�Ę   �������L�D$H�T$H�L$H��hH�L$x�3H  H�D$PH�L$x��G  H�u� H�I`H�L$XH�T$PH�T$HH��$�   H�T$@�D$8    �D$0    �D$(    �D$     E3�D���9   H�D$pH�HH�D$X��  H��h����������L�L$ L�D$H�T$H�L$H��XH�L$h�G  H�D$@H�L$h�?G  H�и H�I`H�L$HH�T$@H�T$0H��$�   H�T$(H��$�   H�T$ L�L$xL�D$p��H�D$`H�HH�D$H���   H��X�������L�L$ L�D$H�T$H�L$H��(H�|$@ tE3��   H�L$8�����H�L$@�H�|$H tE3��   H�L$8�����H�L$H�H�� H�@`L�D$HH�T$@H�L$0H�I���   H��(��������������L�L$ L�D$H�T$H�L$H��(H�ɷ H�@`L�L$HL�D$@H�T$8H�L$0H�I��@  H��(�����������D�D$�T$H�L$H��8�|$P tMH�L$@�͜��H�n� H�I`H�L$ �T$PH��H�D$ ���  H�D$(H�G� H�@`�T$HH�L$(���  �H�+� H�@`�T$HH�L$@H�I���   H��8��������L�L$ L�D$�T$H�L$H��8H�� H�@`H�L$hH�L$(H�L$`H�L$ L�L$XL�D$P�T$HH�L$@H�I���   H��8���������D�L$ D�D$�T$H�L$H��8H��� H�@`�L$h�L$(�L$`�L$ D�L$XD�D$P�T$HH�L$@H�I���   H��8�������������D�L$ D�D$�T$H�L$H��XH�*� H�@`H�D$H    H�D$@    �L$x�L$8��$�   �L$0��$�   �L$(�L$p�L$ E3�D�D$h�3   H�L$`H�I��  H��X����������������������H�T$H�L$H��hH�L$x�D  H��� H�I`H�L$PH�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�D���   H�D$pH�HH�D$P��  H��h�������������������H�T$H�L$H��hH�L$x�xC  H�	� H�I`H�L$PH�D$H    H�D$@    �D$8    �D$0    �D$(    �D$    E3�D���   H�D$pH�HH�D$P��  H��h�������������������H�T$H�L$H��hH�L$x��B  H�y� H�I`H�L$PH�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�D���   H�D$pH�HH�D$P��  H��h�������������������H�T$H�L$H��hH�L$x�B  H�D$PH�L$x�IB  H�ڳ H�I`H�L$XH�T$PH�T$HH�D$@    �D$8    �D$0    �D$(    �D$     E3�D���"   H�D$pH�HH�D$X��  H��h�������������������H�T$H�L$H��hH�L$x��A  H�D$PH�L$x�A  H�:� H�I`H�L$XH�T$PH�T$HH�D$@    �D$8    �D$0    �D$(    �D$     E3�D���5   H�D$pH�HH�D$X��  H��h�������������������D�D$H�T$H�L$H��hH�L$x�SA  H�D$PH�L$x�A  H��� H�I`H�L$XH�T$PH�T$HH�D$@    �D$8    �D$0    �D$(    ��$�   �T$ E3�D���<   H�D$pH�HH�D$X��  H��h�����������L�L$ D�D$�T$H�L$H��XH�
� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �L$p�L$ E3�D�D$h�   H�L$`H�I��  H��� H�@`H�T$xH�L$`H�I���   H��X�������������H�L$H��XH�x� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��   H�L$`H�I��  H��X������������H�T$H�L$H��XH�� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     L�L$hE3��   H�L$`H�I��  H��X���������������������H�L$H��XH��� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��   H�L$`H�I��  H��X�����������̉T$H�L$H��XH�� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�D�D$h�   H�L$`H�I��  H��X����������������������L�D$�T$H�L$H��XH��� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     L�L$pD�D$h�&   H�L$`H�I��  H��X���������������H�L$H��XH�� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��(   H�L$`H�I��  H��X������������H�L$H��XH��� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��#   H�L$`H�I��  H��X������������D�L$ D�D$�T$H�L$H��XH�*� H�@`H�D$H    H�D$@    �D$8    �D$0    �L$x�L$(�L$p�L$ E3�D�D$h�+   H�L$`H�I��  H��X������������H�L$H��hH�L$p����H��� H�I`H�L$PH�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�E3��0   H��H�D$P��  H��h��������������D�D$�T$H�L$H��8H�L$@脒��H�%� H�I`H�L$ �T$HH��H�D$ ��  H��8��������������L�L$ D�D$�T$H�L$H��   H�D$h����H��$�   H�L$p���  �D��$�   �8kdsH�L$p�~���H�D$P    H��$�   ����H��� H�I`H�L$XH�T$PH�T$HH�T$pH�T$@�D$8    ��$�   �T$0��$�   �T$(��$�   �T$ L��$�   D��$�   �2   H��H�D$X��  H�D$PH�D$`H�L$p�y�  H�D$`H�Ę   �������������H�L$H��8H�L$@�=���H�ޫ H�I`H�L$ H��H�D$ ��   H��8����������̉T$H�L$H��XH�D$`H�x u3��YH��� H�@`H�D$H    H�D$@    �D$8    �D$0    �D$(    �D$     E3�D�D$h�-   H�L$`H�I��  H��X����������������������D�L$ L�D$H�T$H�L$H��hL�L$0L�D$<H��$�   H�L$p�|���H�D$LH�D$(H�D$HH�D$ L�L$8L�D$4H�T$xH�L$p������$�    t\��$�    tR�D$49D$<~8�D$H�L$4ȋ�9D$<}&�D$89D$0~�D$L�L$8ȋ�9D$0}
�D$@   ��D$@    �D$@�r�>��$�    t4�D$89D$0~�D$L�L$8ȋ�9D$0}
�D$D   ��D$D    �D$D�2�D$49D$<~�D$H�L$4ȋ�9D$<}
�D$P   ��D$P    �D$PH��h���������������������L�D$H�T$H�L$H��8H�D$PH�D$(H�|$( uH�D$@H��H�D$(E3��diuMH�L$H�H����D$ �|$  u�   �VH�D$(� 9D$ u3��EE3��IicMH�L$H����9D$ uE3��1icMH�L$H�n7  ����t3��H�D$(�L$ ��   H��8���������������L�D$H�T$H�L$H��hH�D$8�����fnicH�L$p�E3  H�D$ H�|$  t�
   H�L$ �Y3  H��t�   A�fnicH�T$@H�L$p�z2  H�D$(H�D$(H�D$0H�T$0H�L$x��  �H�L$@���  H�L$x��3  ���tH�L$x��3  ��u�fnicH�L$x��7  L��$�   �
   H�L$x����H��h����������H�L$H��(H�(� H�@`H�L$0H�I���  H��(���������D�D$H�T$H�L$H��xH�D$8�����mnrsH�L$P���  �D��$�   �   H�L$P����L�L$PL��$�   H�T$@H��$�   �n���H�D$(H�D$(H�D$0H�L$0�E����D$ H�L$@�G����H�L$P���  �D$ H��x��������������������D�D$H�T$H�L$H��xH�D$8������$�    t
�D$ SSSS��D$ DSSS�T$ H�L$P���  �H�L$P�o2  A�   ��H�L$P�����L�L$PL��$�   H�T$@H��$�   螬��H�D$(H�D$(H�D$0H�L$0�u����D$$H�L$@�w����H�L$P��  �D$$H��x��������������������H�L$H��(H�L$0�]���H�D$0H�� H�H�D$0�@   H�D$0�@    H�D$0H��(�������������H�L$H��(H�D$0H�� H�H�L$0�^���H��(����������D�L$ D�D$�T$H�L$H��XH�D$`�@    ��$�    t
�D$@   ��D$@
   �D$8    ��$�   �D$0�D$x�D$(�D$p�D$ D�L$hE3��T$@H�L$`������tH�D$`�x t
�D$D   ��D$D    �D$DH��X��������������̉T$H�L$H��(H�D$0�L$8�HH�L$0荪��H��(���������L�D$H�T$H�L$H��8H�L$H�s0  �D$ �|$ cksat`�|$ TCAbt}�|$ ckhct�|$ atnit��   3���   H�D$@�x t$H�L$@������tH�D$@�@    �   ��   3���   H�D$@�x tH�D$@H� H�L$@�P(�   3��   E3��diemH�L$H�����D$$H�D$@�@   H�D$@H� L�D$H�T$$H�L$@�P �D$,H�D$@�x t�|$$t�|$$u'�|$$u
�D$(   ��D$(    �T$(H�L$@�����D$,�L�D$PH�T$HH�L$@�E���H��8�����������������D�L$ D�D$�T$H�L$H��HH�D$P�x u�1  �D$`�D$ �|$ ��   HcD$ H�
������A H����D$p9D$h~��   �   �D$p9D$h|��   �   �D$p9D$h}��   �   �D$p9D$h�   �r�D$p9D$h~�D$x9D$h}�   �W�D$p9D$h|�D$x9D$h�   �<�D$p9D$h|�D$x9D$h}�m�$�D$p9D$h~�D$x9D$h�U��D$p9D$ht�G�T$XH�L$(��#  H�T$(H�L$P�����*D$x�*L$pA�   (ЋL$`�d�  H�D$P�@    H��H� @ @ *@ >@ O@ j@ �@ �@ �@ �������������\$ D�D$�T$H�L$H��HH�D$P�x u�i  �D$`�D$ �|$ �  HcD$ H�y�������B H����D$hf/D$pv�+  ��   �D$hf/D$pr�  ��   �D$pf/D$hv��   �   �D$pf/D$hr��   �   �D$hf/D$pv�D$xf/D$hv�   �u�D$hf/D$pr�D$xf/D$hr�   �R�D$hf/D$pr�D$xf/D$hv�z�2�D$hf/D$pv�D$xf/D$hr�Z��D$hf.D$pzt�F�T$XH�L$(�"  H�T$(H�L$P�8���D��$�   �T$x�L$p�L$`��  H�D$P�@    H��H�f��A �A �A �A �A B 9B YB yB ���������������������\$ D�D$�T$H�L$H��H�D$0   �D$x�D$(�D$p�D$ �\$hD�D$`�T$XH�L$P�����H��H������������\$ D�D$�T$H�L$H��H�D$0   �D$x�D$(�D$p�D$ �\$hD�D$`�T$XH�L$P����H��H������������\$ D�D$�T$H�L$H��H�D$0   �D$x�D$(�D$p�D$ �\$hD�D$`�T$XH�L$P����H��H�����������H�L$H��(H�L$0����H�D$0H��� H�H�D$0�@   H�D$0H��(���������H�L$H��(H�D$0H��� H�H�L$0�.���H��(����������L�D$H�T$H�L$H��8H�L$H�#*  �D$ �|$ cksat=�|$ ckhct�RH�D$@�@   H�L$@�S�����tH�D$@�@    �   �93��5H�D$@�x tH�D$@H� H�L$@�P(�3��L�D$PH�T$HH�L$@裠��H��8���������������L�D$H�T$H�L$H��8H�D$ ����H�L$@�����H�D$@H�� H�H�D$@H�L$PH�H(E3��myalH�L$H����H�L$@�A H�D$@�x tH�D$@�x tH�D$@�@     A�
   �hfedH�L$H�H���H�L$@�A$H�D$@H��8����������L�D$H�T$H�L$H��8H�L$H��(  �D$ �|$ ytsdt�!H�L$@�I���H�D$@H� H�L$@�P8�   �L�D$PH�T$HH�L$@�>���H��8����������H�L$3����������H�L$3����������H�L$�����������H�L$3����������H�L$3����������H�L$3����������H�T$H�L$3���������������������H�T$H�L$H��XH�D$(�����D$     H�L$0��  �H�T$0H�L$h�  �D$ ���D$ H�L$0�r  H�D$hH��X���������H�L$H��H�D$ H�x( u3��%H�D$ H�@(� ����t	�$   ��$    �$H����������������H�L$����������̉T$H�L$H��(H�D$0H� H�L$0���   ��t-H�D$0�L$89H tH�D$0�L$8�H H�D$0H� H�L$0���   H��(�����������H�L$H�D$�@ �������������������H�L$H��(�0   3��  ��H�L$0�O�  H��(����������̉L$H��8�0   3��  �D$ �L$@�?����L$ ��H����  H��8�������������H�T$�L$H��hH�D$8�����0   3��>  �D$ L�D$x�T$pH�L$@����H�D$(H�D$(H�D$0�D$ ��H�L$0��  �H�L$@�����H��h���������L�D$H�T$�L$H��hH�D$8�����0   3���  �D$ L��$�   L�D$x�T$pH�L$@�����H�D$(H�D$(H�D$0�D$ ��H�L$0�+�  �H�L$@�k���H��h������������H�L$H��8�    �   �X  ��H�L$@���  ��u
�D$    ��D$     �D$ H��8������������̉L$H��8�    �   �	  �D$$�L$@�����L$$��H����  ��u
�D$    ��D$     �D$ H��8���������������H�T$�L$H��hH�D$@�����    �   �  �D$$L�D$x�T$pH�L$H�t���H�D$0H�D$0H�D$8�D$$��H�L$8��  ��u
�D$    ��D$     �D$ �D$(H�L$H�'����D$(H��h��������������������L�D$H�T$�L$H��hH�D$@�����    �   ��  �D$$L��$�   L�D$x�T$pH�L$H����H�D$0H�D$0H�D$8�D$$��H�L$8�X�  ��u
�D$    ��D$     �D$ �D$(H�L$H�z����D$(H��h�������H�T$�L$H��(H�� H�@L�D$8�T$03����  H��(�������������������L�D$�T$�L$H��(H��� H�@L�L$@D�D$8�T$03����  H��(����������L�L$ D�D$�T$H�L$H��8H�Z� H�@H�L$hH�L$(�L$`�L$ L�L$XD�D$P�T$HH�L$@���  H��8���������������H�L$H��(H�� H�@`H�L$0���  H��(�������������D�D$�T$H�L$H��hH�D$8�����D$     H��� H�@`D��$�   �T$xH�L$@���  H�D$(H�D$(H�D$0H�T$0H�L$p�����D$ ���D$ H�L$@�����H�D$pH��h���������������H�T$H�L$H��   H�D$p�����D$(    H�L$@�"�����D$     �
�D$ ���D$ 3�����   �D$ k�
E3���H��$�   �����D$,�D$ k�
��E3���H��$�   �����D$$�|$$ u�w�|$  ~/E3�H�2� H�L$X�����H�T$XH�L$@�D  �H�L$X����D�D$$�T$,H�L$x����H�D$0H�D$0H�D$8H�T$8H�L$@�  �H�L$x������/���H�T$@H��$�   �f����D$(���D$(H�L$@����H��$�   H�Ę   ������������������H�T$H�L$H��(H�� H�@`H�T$8H�L$0���  H��(�������������������D�L$ D�D$�T$�L$H��8H��� H�@`H�L$hH�L$(�L$`�L$ D�L$XD�D$P�T$H�L$@���  H��8����������������̉L$H��(H�Y� H�@`�L$0���  H��(���������������H�L$H��(W�H�D$0H�H�	  H�D$0H�@H�L$0H�IH� H�T$0�PHE3�3ҹ�����  H��(����������������������H�L$H�D� ��������������������H�L$H��h  HǄ$�   ����H��$p  H� H��$(  H��$p  �PPH��$�   H��$�   H��$�   H��$�   H��$p  �͛���H��$(  ����H��$�   �0���H�D$xH�D$xH��$�   �D$@    �D$8    �D$0    H��$�   H�D$(�D$     A�   A�?   3�H��$p  ������H��$�   �E���H��$�   軿��H��$�   H��$�   H��$�   �(   ��"  �D$0    H��$�   H�L$(�D$     D��A�   ��  H��$p  �����H��u
�D$T   ��D$T    �D$T�D$PH��$�   豿���D$P��t3��  H��$�   ����H��$�   H��$�   H�D$`�D$@    �D$8    �D$0    H�D$`H�D$(�D$     E3�A�8   3�H��$p  ������H��$�   �/����   H��$p  �R���H��$@  �E�  H��$�   H��$�   H�D$p�   ��!  �D$X�,  �!  �D$\H��$  �U���H�D$hH�D$hH��$�   H�D$pH�D$8�D$X�D$0�D$\�D$(�D$ ;   L��$�   A�	����  H��$p  �����H��$  �p����H��$@  �W�  H��$p  ����H��$p  �����   H��$p  �{���H��$p  H��$p  H�H8�   ��  �   H��h  �����������������H�L$H��hH�D$0����H�D$pH�� �   H���8�  H�D$pH�@P    H�D$pH�@X    H�D$pH�@`    H�D$pW��@@��   H�L$p�U���E3�H��� H�L$H�m������  H�L$8�1  �D$     E3�L�D$HH�T$8H�L$p�¢���H�L$H�B���H�D$pH�� E3��   H���.�  H��h����������H�T$H�L$H���   H�D$x����E3�H�T� H��$�   �ۼ�����  H�L$h�  H��$   �@@�Y� �,���H��$�   輼��H�D$@H�D$@H�D$8L��$�   H�T$8H��$�   �  H�D$0H�D$0H�D$H�D$     E3�L�D$HH�T$hH��$   �͡���H��$�   �J����H��$�   �<����H��$�   �.����tatsH�L$P蔼  �A�   �   H�L$P�n  H��$   �P@�   H�L$P�B  ��  H��$�   �  L�L$PL��$�   H��$�   H��$   ����H��$�   �n��H��$   H�xP ��   H��$   H��HH���  H��$   H�xP tEH��$   H�HXH��$   �PPH��$   H�A`H��$   H�@X    H��$   H�@P    �H��� ��  �u��H��$   H��HH���Q  �H�L$P���  H���   ���������������L�D$H�T$H�L$H��   H�D$P����H��$�   �  �D$ �|$ MicM��   �|$ ckhctq�|$ fnict�+  �   H�L$x���  H�D$(H�D$(H�D$0H�T$0H��$�   �y�  �H�L$x�N�  A�   �   H��$�   衹���   ��   ��   H��$�   H� H��$�   �P(��u3���   �   �   �   E3��IicMH��$�   �/����D$$�|$$���t�t�tatsH�L$8�C�  �E3��   H�L$8�   ��  H�L$X�q  L�L$8L�D$XH�T$hH��$�   ����H�L$h��k���H�L$8�p�  �   H��$�   ����L��$�   H��$�   H��$�   ����H�Ę   ����������L�D$�T$H�L$H��8�D$H�D$ �|$ t�3H�D$@H�� �   H���g�  �   �}�  3�H�L$@�!����   �L�D$P�T$HH�L$@�g���H��8�������������������H�L$H��(H�D$0H�� �   H����  �   ��  3�H��(������������������L$H�L$H�D$�D$�@@���������������������H�L$H�D$H�� ������������������L�D$H�T$H�L$H��8H�D$     3����,  H�D$@H�xP t9H�� �~  ��q���
   �b�  H�D$@H�� H����  ��t3���   �H�D$@H��HH���  H�D$@H�xP ��   H�D$@H�L$PH�HXH�D$@H�L$HH�HPH�D$@H��HH���  H�D$@H�xP t%�
   ���  H�D$@H�� H���_  ��t3��o��H�D$@H��HH���4  H�D$@H�@`H�D$ H�D$@H�@`    H�D$@H��HH���H  �)�"H�5� ��  ��p��H�D$@H��HH���"  �����H�D$ H��8��������������������L�D$H�T$H�L$H��hH�D$X�����D$     H�L$@�¶  �H�|$x t^H�
� H�@hH�L$x�PH�D$(H�|$( u�D$8    H�L$@�G�  �D$8�   H�D$(H� L�D$@H��$�   H�L$(�PP�D$ �YH��� H�@`H�L$p�PH�D$0H�|$0 u�D$<    H�L$@��  �D$<�aH�D$0H� L�D$@H��$�   H�L$0�P@�D$ H�L$@�  ���tH�D� H�@`H�T$@H�L$p���   �D$ �D$$H�L$@膶  �D$$H��h��������������D�D$H�T$H�L$H��8E3��T$PH�L$H虴���D$ �T$ H�L$@�  H��8����������������������D�L$ L�D$H�T$H�L$H��H�D$p9D$hu,E3��tsemH�L$`�9�����uE3��rdemH�L$`�#�����t3��E�D$     �T$hH�L$(�  L�D$ H�T$(H�L$X������u3���T$ H�L$P��  �   H��H���������������������D�D$H�T$H�L$H���   H�D$h����H�L$P�ճ���H�L$p�ʳ��H�D$(H�D$(H�D$HL�L$HD��$�   H��$�   H��$�   �;���H�D$@H�D$@H�D$8H�T$8H�L$P�=+���H��$�   �����H�L$p�߳��H��$�   H�D$0H�T$PH�L$0�x���H�D$ H�T$ H��$�   ��  �H�L$P衳��H���   ���������������D�L$ L�D$H�T$H�L$H��   H�D$`������$�   9�$�   u2E3��tsemH��$�   脲����uE3��rdemH��$�   �k�����t3��   H�L$8藲�����$�   H�L$P��  L�D$8H�T$PH��$�   谜����u�D$     H�L$8�ղ���D$ �FH�D$hH�D$0H�T$8H�L$0�k���H�D$(H�T$(H��$�   ��  �D$$   H�L$8荲���D$$H�Ĉ   �������D�D$H�T$H�L$H��8E3��T$PH�L$H�l  �D$ �T$ H�L$@�J  H��8����������������������D�L$ L�D$H�T$H�L$H��H�D$p9D$hu,E3��tsemH�L$`�9�����uE3��rdemH�L$`�#�����t3��E�D$     �T$hH�L$(�  L�D$ H�T$(H�L$X�4�����u3���T$ H�L$P�
  �   H��H���������������������D�D$H�T$H�L$H��8WҋT$PH�L$H�  �D$ �L$ H�L$@�  H��8������������������D�L$ L�D$H�T$H�L$H��H�D$p9D$hu,E3��tsemH�L$`�9�����uE3��rdemH�L$`�#�����t3��HW��D$ �T$hH�L$(�  L�D$ H�T$(H�L$X�c�����u3���L$ H�L$P�[
  �   H��H������������������D�D$H�T$H�L$VWH��   H�L$ �6���H�L$`�,���L��D��$�   H�T$xH��$�   胯��H�L$ H��H��   �H�D$@H�L$ H��H��   �H�T$@H��$�   �
  H�Ę   _^�������������������D�L$ L�D$H�T$H�L$VWH��   ��$�   9�$�   t'��$�   9�$�   t��$�   9�$�   t3���   E3��tsemH��$�   贮����uE3��rdemH��$�   蛮����t3��   W�H�L$`��  ��$�   H�L$0��  ��$�   H�L$@��  ��$�   H�L$P��  H�D$`H�D$ L�L$0L�D$@H�T$PH��$�   ������u3��4H��$�   H�L$`H��H��   �H��$�   H��$�   ��  �   H�Ĩ   _^��������D�D$H�T$H�L$VWH��hH�L$ �  H�L$@�  L��D��$�   H�T$PH��$�   ��  H�L$ H��H��   �H�D$0H�L$ H��H��   �H�T$0H��$�   �  H��h_^���������L�L$ L�D$H�T$H�L$VWH��X��$�   9�$�   u2E3��tsemH��$�   ������uE3��rdemH��$�   �������t3��jH�L$ �6  ��$�   H�L$0�U  L�L$ L��$�   H�T$0H�L$x�ɘ����u3��+H�D$@H�L$ H��H��   �H�T$@H�L$p��  �   H��X_^����������������H�T$H�L$H��(H�D$0H�L$8�	�H�D$8H��H�L$0H��H���J^��H�D$0H��(�H�L$H��XH�D$0����H�D$`H��H���  �H�D$`� ����H�L$8�  H�D$ H�D$ H�D$(H�D$`H��H�T$(H���  �H�L$8��^���H�D$`H��X�������������H�L$H�D$W�� H�D$��� �@H�D$�������̉T$H�L$H�D$�L$�H�D$H�@    H�D$���������̉T$H�L$H�D$�    H�D$�L$�HH�D$����������̉T$H�L$H�D$�    H�D$�L$�HH�D$�����������H�L$H�D$�     H�D$�@    H�D$����������������L$H�L$H�D$�D$� H�D$�D$�@H�D$�D$�@H�D$�H�L$H��(H�D$0H��H���v]��H��(��H�L$H��(H�L$0����H��(���������H�T$H�L$H��(E3�H�T$0H�L$8�  H�D$0H��(�������H�T$H�L$H��H�D$ H�L$(� f.z;u9H�D$ H�L$(�@f.Az#u!H�D$ H�L$(�@f.Azu	�$    ��$   �$H�������H�T$H�L$H��8H�D$@H�L$H� f.zuH�D$@H�L$H�@f.Azu3��]H�D$@H�L$H� �YA��  �D$(H�D$HH�L$@��YI(���  �L$(f.�zt
�D$    ��D$     �D$ H��8���������������H�T$H�L$H��8H�T$HH�L$@������t
�D$    ��D$     �D$ H��8�����L�D$H�T$H�L$H��XH�D$(�����D$     H�T$hH�L$0�����H�T$pH�L$0�]   H�T$0H�L$`�Ψ���D$ ���D$ H�L$0����H�D$`H��X���������������̉T$�L$�D$�L$ȋ�������������H�T$H�L$H��8H�L$@��  �D$ ����A�����L�D$H��H�L$@����H�D$@H��8���������������̉T$H�L$H��(H�L$0�9|���D$8����t
H�L$0�J���H�D$0H��(����������̉T$H�L$H��(H�L$0�y����D$8����t
H�L$0�
���H�D$0H��(����������̉T$H�L$H��(H�L$0�Yb���D$8����t
H�L$0�ʧ��H�D$0H��(����������̉T$H�L$H��(H�L$0褧���D$8����t
H�L$0芧��H�D$0H��(����������̉T$H�L$H��(H�L$0������D$8����t
H�L$0�J���H�D$0H��(����������̉T$H�L$H��(H�L$0�	����D$8����t
H�L$0�
���H�D$0H��(����������̉T$H�L$H�D$�8�uH�D$�     H�D$�L$�H�#H�D$�8 uH�D$�L$9HtH�D$�    ����������������̉T$H�L$H�D$�8�uH�D$�     H�D$�L$�H�#H�D$�8 uH�D$�L$9HtH�D$�    ������������������L$H�L$H�D$�8�uH�D$�     H�D$�D$�@�)H�D$�8 uH�D$�@f.D$ztH�D$�    �����H�T$H�L$VWH��(H�D$@�8�u"H�D$@�     H�D$@H�xH�t$H�   ��/H�D$@�8 u%H�D$@H��H�T$HH��������tH�D$@�    H��(_^���������������H�T$H�L$VWH��(H�D$@�8�u"H�D$@�     H�D$@H�xH�t$H�   ��/H�D$@�8 u%H�D$@H��H�T$HH��������tH�D$@�    H��(_^���������������H�T$H�L$H��8H�D$ ����H�D$@�8�u#H�D$@�     H�D$@H��H�T$HH�������/H�D$@�8 u%H�D$@H��H�T$HH���������tH�D$@�    H�L$H�^���H��8���������������L�D$H�T$H�L$H��(H��v H��  L�D$@H�T$0H�L$8�PH��(����������D$H��(�D$0�z� H��(������D�D$�T$H�L$H��(H�_v H�@ D�D$@�T$8H�L$0��8  H��(�����������D�D$H�T$H�L$H��hH�D$8�����D$     H�v H�@ D��$�   H�T$@H�L$p���   H�D$(H�D$(H�D$0H�T$0H�L$x���  �D$ ���D$ H�L$@�&�  H�D$xH��h������������̉T$H�L$H��(H��u H�@ �T$8H�L$0���   H��(����̉T$H�L$H��(H�du H�@ �T$8H�L$0���  H��(�����H�L$H�D$�@�L�L$ D�D$H�T$H�L$H��xH�D$8�����D$     H�u H�@ L��$�   D��$�   H�T$@H��$�   ��P  H�D$(H�D$(H�D$0H�T$0H��$�   �����D$ ���D$ H�L$@�s���H��$�   H��x�������H�L$H��(H��t H�@ H�L$0�P@H��(����������������H�L$H��(H�Xt H�@(H�L$0�PxH��(����������������H�L$H�D$� ���T$�T$H�L$H��(H�t H�@ �T$@�T$8H�L$0��0  H��(���������L�L$ D�D$H�T$H�L$VWH��8H��s H�@ L�L$hD�D$`H�T$ H�L$P��X  H�|$XH��   �H�D$XH��8_^�������H�L$H��H�D$ �8u	�$   ��$    �$H��������H�L$H��H�D$ �8u	�$   ��$    �$H��������H�L$H��H�D$ �8u	�$   ��$    �$H��������H�L$H��H�D$ �8u	�$   ��$    �$H��������H�L$H��H�D$ �8u	�$   ��$    �$H��������H�L$H��(H��r H��  H�L$0�PH��(�������������H�L$H�D$H����H�L$H�D$H����H�L$H�D$H����H�L$H�D$H����H�L$H�D$H����H�L$H�D$H����H�L$H��(H��q H��  H�L$0���   H��(����������L�D$�T$H�L$H��(H��q H�@ L�D$@�T$8H�L$0��x  H��(�����������H�L$H�D$� ����H�L$H��(H�xq H���   H�L$0���   H��(����������H�L$H�D$H�@���D$�D$�Y�� �^�� ����D�D$�T$H�L$H��(H�q H�@ D�D$@�T$8H�L$0�P`H��(��������������L�D$�T$H�L$H��(H��p H�@ L�D$@�T$8H�L$0��  H��(�����������L�D$�T$H�L$H��(H��p H�@ L�D$@�T$8H�L$0�PxH��(�������������̉T$H�L$H��(H�Tp H�@ �T$8H�L$0�PHH��(���������T$�T$H�L$H��(H�p H�@ �T$@�T$8H�L$0�PXH��(������������L�D$�T$H�L$H��(H��o H�@ L�D$@�T$8H�L$0���   H��(����������̉L$H��(3ҋL$0�   H��(��������̉T$�L$�D$��D$�������������H�L$H��(H�ho H���   H�L$0H�I�P(H��(���������H�L$H��(H�8o H���   H�L$0���   H��(�����������L$H�L$H��(H�o H���   �L$8H�L$0�PH��(�����������������H�L$H��(H��n H���   3�H�L$0��  H��(�������̉T$H�L$H��(H��n H���   D�D$83�H�L$0��  H��(���������������H�L$H��(H�Xn H���   �   H�L$0��  H��(��������������������̉T$H�L$H��(H�n H���   D�D$8�   H�L$0��  H��(������������H�L$H��8H��m H���   �   H�L$@��  ��t
�D$    ��D$     �D$ H��8����������̉T$H�L$H��(H��m H���   D�D$8�   H�L$0��  H��(������������H�L$H��(H�Hm H���   H�L$0���  H��(���������̉T$H�L$H��(H�m H���   �T$8H�L$0���  H��(������������������H�T$H�L$H��(H��l H���   H�T$8H�L$0���  H��(���������������̉T$H�L$H��(H��l H���   �T$8H�L$0���  H��(������������������D�D$�T$H�L$H��(H�Ol H���   D�D$@�T$8H�L$0��0  H��(��������D�D$H�T$H�L$H��(H�l H���   D�D$@H�T$8H�L$0��8  H��(����������������������H�L$H��(H��k H���   H�L$0��   H��(����������L�D$�T$H�L$H��8�L$H�5 H�D$ H�|$  tL�D$PH�T$ H�L$@�t   H�D$ H��8�����������L�L$ D�D$�T$H�L$H��8�T$P�L$H� H�D$ H�|$  tL�D$XH�T$ H�L$@�   H�D$ H��8������������������L�D$H�T$H�L$H��(H��j H���   L�D$@H�T$8H�L$0��@  H��(����������������������D�D$�T$H�L$H��(H��j H���   D�D$@�T$8H�L$0��H  H��(��������H�T$H�L$H��(H�Sj H���   H�T$8H�L$0���  H��(����������������H�L$H��(H�j H���   H�L$0��x  H��(����������D�L$ D�D$H�T$H�L$H��8H��i H���   H�L$hH�L$(�L$`�L$ D�L$XD�D$PH�T$HH�L$@��h  H��8�����������\$ D�D$�T$H�L$H��XH�D$0����E3���  H�L$`�����|$h u�   �E3���  H�L$`����H�D$(H�|$( u3��\H�L$8�Җ  �D�D$p��  H�L$8������T$x��  H�L$8�����E3�H�T$8H�L$(��G  �D$    H�L$8�D�  �D$ H��X������������H�L$H��(H��h H���   H�L$0���  H��(����������H�T$H�L$H��(H��h H���   H�T$8H�L$0��`  H��(����������������H�T$H�L$H��(H�Ch H���   H�T$8H�L$0��X  H��(����������������H�L$H��(H�h H���   H�L$0��h  H��(���������̉L$H��(H��g H���   �L$0�H��(����������������H�L$H��(H��g H���   H�L$0H�	�P H�D$0H�     H��(��������������D�L$ L�D$H�T$H�L$H��XH�D$@    H�D$8    H�D$H    H��$�   �8 u0H�T$hH�L$`�9  ��u�   H�L$`�~C  ��u
�D$0    ��D$0   H��$�   �L$0�H��$�   �8 ��   H�L$`�_  ��$�    u5H��$�   H�D$(H��$�   H�D$ D�L$xL�D$pH�T$hH�L$`��  �XH�D$pH�D$8�H�L$8�z=  H�D$8H�|$8 t5H��$�   H�D$(H��$�   H�D$ D�L$xL�D$8H�T$hH�L$`�j  �H��$�   �8 uH�L$`��  ��t
�D$4    ��D$4   H��$�   �L$4�H��$�   �8 uH�L$`�&  H�T$hH�L$`�;  ��   H�L$`�X  ��$�    u9H��$�   H�D$(H�D$     D�L$xL�D$pH�T$hH�L$`�   H�D$@�   �  ����H�D$@H�|$@ u3��   H�L$p�-<  H��H�L$@�D  H�D$pH�D$8�H�L$8�:<  H�D$8H�|$8 tMH��$�   H�D$(H�D$     D�L$xL�D$8H�T$hH�L$`�.   H�D$HH�|$H tH�T$@H�L$H�>  �H�D$@H��X�������D�L$ L�D$H�T$H�L$H��8H��d H���   H�L$hH�L$(H�L$`H�L$ D�L$XL�D$PH�T$HH�L$@��p  H��8��������H�L$H��(H�hd H���   H�L$0���  H��(����������H�L$H��(H�8d H���   H�L$0���  H��(����������L�D$H�T$H�L$H��(H��c H���   L�D$@H�T$8H�L$0���  H��(����������������������H�L$H��(H��c H���   H�L$0���  H��(����������H�L$H��(H��c H���   H�L$0���  H��(����������H�L$H��(H�Xc H���   H�L$0���  H��(����������H�L$H��(H�(c H���   H�L$0���  H��(����������H�L$H��(H��b H���   H�L$0���  H��(����������H�T$H�L$VWH��HH��b H���   H�T$`H�L$ ���  H�|$hH��   �H�D$hH��H_^��������H�L$H��(H�xb H���   H�L$0���  H��(���������̉T$H�L$H��(H�Db H���   �T$8H�L$0���  H��(�������������������L$H�L$H��(H�b H���   �L$8H�L$0���  H��(���������������L$H�L$H��(H��a H���   �L$8H�L$0���  H��(���������������L$H�L$H��(H��a H���   �L$8H�L$0���  H��(��������������H�T$H�L$H��(H�Ca H���   H�T$8H�L$0���  H��(����������������L�L$ L�D$H�T$H�L$H��8H��` H���   �L$`�L$ L�L$XL�D$PH�T$HH�L$@��  H��8��������������������L�L$ L�D$H�T$H�L$H��HH��` H���   ��$�   �L$0H�L$xH�L$(�L$p�L$ L�L$hL�D$`H�T$XH�L$P��  H��H���������������H��(H�=` H���   ��  �H��(�������������������H�L$H��(H�` H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H��_ H���   H�L$0���  H��(����������H�L$H��(H��_ H���   H�L$0���  H��(����������H�T$H�L$H��(H�c_ H���   H�T$8H�L$0���  H��(���������������̉T$H�L$H��(H�$_ H���   �T$8H�L$0���  H��(������������������L�D$�T$H�L$H��(H��^ H���   L�D$@�T$8H�L$0��@  H��(��������D�D$�T$H�L$H��(H��^ H���   D�D$@�T$8H�L$0��   H��(��������L�D$�L$H�L$H��(H�]^ H���   L�D$@�L$8H�L$0��  H��(�������������������̉T$�L$H��8�  �*���H�D$ H�|$  u3��   E3�D�D$@��  H�L$ ����H��u�;�9E3�D�D$H�(  H�L$ �o���H��u��E3��   H�L$ �d<  H�D$ �)H�|$  tH��] H���   H�L$ �P H�D$     3�H��8����������������H�L$H��(H�X] H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H�] H���   H�L$0��  H��(����������H�L$H��(H��\ H���   H�L$0��  H��(����������H�L$H��(H��\ H���   H�L$0��H  H��(����������H�L$H��(H��\ H���   H�L$0��P  H��(����������H�L$H��(H�X\ H���   H�L$0���  H��(����������D�D$�T$H�L$H��(H�\ H���   D�D$@�T$8H�L$0��  H��(��������D�L$ D�D$�T$H�L$H��(H��[ H���   D�L$HD�D$@�T$8H�L$0��   H��(��������������D�L$ D�D$�T$H�L$H��8H��[ H���   �L$`�L$ D�L$XD�D$P�T$HH�L$@���  H��8����������������������D�D$H�T$H�L$H��8H�D$     �|$PuH�L$@����H�D$ �.�|$P uH�L$@�;���H�D$ ��|$PuH�L$@����H�D$ H�|$  u3��L�D$ H�T$HH�L$@�   H��8����������L�D$H�T$H�L$H��h�� H�D$HH�|$H tH��$�    u3��-  H�L$p�/2  H�D$PH�L$p� 2  ���D$<H�|$P u
H�D$H��   �D$4    �
�D$4���D$4H��$�   �V
 9D$4��   H�D$DH�D$ L�L$@D�D$<�T$4H��$�   �� ��u봋D$@�D$0�
�D$0���D$0�D$D9D$0}�D$0����u2�D$0��H�Hk��L$0��Hc�Hk�H�T$PL�D$PA�L9Lu뮋D$0����H�L$x��0  �L$0��HcɋD��D$8�|$8�t�T$8H�L$H�	 �o�������H�D$HH��h��������D�L$ L�D$H�T$H�L$H��HH�L$P��0  H�D$8H�|$8 u3��  H�D$(    �|$huH�L$P�`���H�D$(�.�|$h uH�L$P����H�D$(��|$huH�L$P�`���H�D$(H�|$( u3��X  H�L$(��	 �D$     �
�D$ ���D$ H�L$P�$0  9D$ �!  �T$ H�L$X��/  H�D$0H�|$0 u�Ÿ   Hk� H�L$0�TH�L$`�Q5  ��t�D$ ����H�L$(� �   Hk�H�L$0�TH�L$`�5  ��t�D$ ��   ��H�L$(�S HcD$ Hk�HcL$ Hk�H�T$8L�D$8A�L9Lt7�   Hk�H�L$0�TH�L$`��4  ��t�D$ ��   ��H�L$(�� �   Hk�H�L$0�TH�L$`�4  ��t�D$ ��   ��H�L$(� ������   H��H����������������H�L$H��(H�8W H���   H�L$0���  H��(����������L�D$H�T$H�L$H��(H��V H���   L�D$@H�T$8H�L$0���  H��(����������������������L�L$ L�D$�T$H�L$H��(H��V H���   L�L$HL�D$@�T$8H�L$0���  H��(��������������H�L$H��(H�hV H���   H�L$0���  H��(����������H�L$H��(H�8V H���   H�L$0���  H��(����������H�T$H�L$H��(H�V H���   H�T$8H�L$0��  H��(����������������H�T$H�L$H��(H��U H���   H�T$8H�L$0��  H��(����������������H�L$H��(H��U H���   H�L$0��  H��(����������H�T$H�L$H��(H�SU H���   H�T$8H�L$0��   H��(����������������H�L$H��(H�U H���   H�L$0���  H��(����������D�D$H�T$H�L$H��(H��T H���   D�D$@H�T$8H�L$0��(  H��(����������������������H�T$H�L$H��(H��T H���   H�T$8H�L$0��p  H��(����������������H�T$H�L$H��(H�ST H���   H�T$8H�L$0��x  H��(����������������D�L$ D�D$H�T$H�L$H��(H�	T H���   D�L$HD�D$@H�T$8H�L$0���  H��(�����������̉T$H�L$H��(H��S H���   �T$8H�L$0��(  H��(������������������H�T$H�L$H��(H��S H���   H�T$8H�L$0���  H��(����������������H�L$H��(H�HS H���   H�L$0���  H��(���������̉T$�L$H��8��  �*���H�D$ H�|$  u3��CD�D$H�T$@H�L$ ������u'H�|$  tH��R H���   H�L$ �P H�D$     H�D$ H��8������������������H�L$H��(H��R H���   H�L$0H�	�P H�D$0H�     H��(��������������L�L$ D�D$H�T$H�L$H��(H�IR H���   L�L$HD�D$@H�T$8H�L$0��@  H��(�������������L$H�L$H��(H�R H���   �L$8H�L$0��H  H��(��������������H�L$H��(H��Q H���   H�L$0��P  H��(����������D�D$�T$H�L$H��(H��Q H���   D�D$@�T$8H�L$0��X  H��(��������H��(H�]Q H���   ��0  H��(��������������������H�L$H��(H�(Q H���   H�L$0��8  H��(����������H�L$H��8H�L$@��&  E3���  H���}���D$ H�L$@��'  ���|$ u�D$ ��3�H��8���������������������H�L$H��(H�L$0��}��E3���  H������H��(���������D�L$ �T$H�T$H�L$VWH��XH�VP H���   H��$�   H�L$ D��$�   ��$�   H�T$pH�L$0��   H�|$xH��   �H�D$xH��X_^���������������D�L$ �T$H�T$H�L$VWH��XH��O H���   H��$�   H�L$ D��$�   ��$�   H�T$pH�L$0��(  H�|$xH��   �H�D$xH��X_^���������������H�L$H��(H�hO H���   H�L$0��8  H��(����������D�D$�T$H�L$H��(H�/O H���   D�D$@�T$8H�L$0��p  H��(��������L�L$ �T$H�T$H�L$H��(H��N H���   L�L$H�T$@H�T$8H�L$0��`  H��(���������̉T$�L$H��(H��N H���   �T$8�L$0�PH��(�������H�L$H��(H�xN H���   H�L$0H�	�P H�D$0H�     H��(���������������\$ L�D$�T$H�L$H��8H�)N H���   H�L$hH�L$(�L$`�L$ �\$XL�D$P�T$HH�L$@���  H��8�����������\$ L�D$�T$H�L$H��8H��M H���   H�L$`H�L$ �\$XL�D$P�T$HH�L$@���  H��8������������������H�L$H�D$H�     H�D$����������H�L$H��(H�XM H���   �   H�L$0H�	���  H��(������������������H�T$H�L$H��8H�M H���   H�L$H���  H�L$@H�H�D$@H�8 t
�D$    ��D$     �D$ H��8������������H�L$H��(H��L H���   3�H�L$0H�	���  H��(���������������������D�L$ D�D$�L$�L$H��(�*D$0�YD$8�X� �,��D$0D�D$H�T$@�L$0�z)  H��(����������������������H�L$VWH��  H��$�  �5#  �D$D�D$$    H��$�  �<#  H�D$hH�D$x    H�D$H    HǄ$�       H�D$X    �|$D u
�   �  H��$�  ��$  =�  ��  E3��:  H��$�  ��#  H��$�   H��$�  �#  ��$�   Ǆ$�       H��$�  �.#  H�D$8H��$�  ����H��$�   H��$�  ����H��$�   �D$     �
�D$ ���D$ ��$�   9D$ �  H��$�    ��   A������T$ H��$�   ��  �D$@�|$@���   HcD$@Hk�H��$�   H�H��H���&!  9D$ t�HcD$@Hk�H��$�   H�H��H���/ ��$�   ��$�   9�$�   ~��$�   ��$�   HcD$@Hk�H��$�   H�H��H���{ �L$$ȋ��D$$�?HcD$ Hk�HcL$ Hk�H�T$8L�D$8A�L9Lu�D$$���D$$��D$$���D$$�����H��$�    t&E3�H��$�  H��$�   �F�  ��u
�  �  H��$�    ��   H��$�   ��  H����   H��$�   ��  ;D$DunHcD$DHk�H�xI H�IH��$`  L�]� ��  ��H��$`  ��P  H�D$xH�|$x u
�  ��  H��$�   �D�  D�D$DH�T$xH���  HcD$DHk�H�
I H�IH��$   L�� ��  ��H��$   ��P  H�D$HH�|$H u
�  �  D�D$DH�T$HH�L$h�  ��$�    ~V��$�   ��H�H��H��H H�IH��$@  L�˥ ��  ��H��$@  ���  H�D$XH�|$X u
�!  �  A������T$$H��$�  ������u
��  ��  H��$�    t)A�   H��$�  H��$�   ��  ��u
��  ��  H��$�    tH��$�   �.�  H��$�   �HǄ$�       H��$�   H��$�   H��$�  ��  H�D$h�D$$    �D$     �
�D$ ���D$ ��$�   9D$ �t  H��$�    ��  A������T$ H��$�   �s �D$@�|$@���  HcD$@Hk�H��$�   H�H��H���  9D$ t�HcD$@Hk�H��$�   H�H��H���> ��$�   �D$p    �D$(    �D$t    �
�D$t���D$tHcD$@Hk�H��$�   H�H��H���  9D$t��  HcD$@Hk�H��$�   H�H���T$tH���'#  ��u�HcD$@Hk�H��$�   H�H���T$tH���  �D$0HcD$0Hk�HcL$(H�T$XL�D$8A� ���D$(���D$(�D$0��HcL$(H�T$X���D$(���D$(HcD$0Hk�HcL$(H�T$XL�D$8A�D ���D$(���D$(�D$0��   HcL$(H�T$X���D$(���D$(HcD$0Hk�HcL$(H�T$XL�D$8A�D ���D$(���D$(�D$0��   HcL$(H�T$X���D$(���D$(HcD$0Hk�HcL$(H�T$XL�D$8A�D ���D$(���D$(�D$0��   HcL$(H�T$X���D$(���D$(�M����D$(��$�   ��$�    ��  ��$�   �+���H�L��H�T$XH��$�   �n  �D$(    ��$�   9D$p|1L�J� A�  H�M� H�n� �9�  H�r� �  �,����$�   9D$p|
�c
  �^
  HcD$(H�L$X����$�   H��$�    t1Hc�$�   Hk�HcL$$Hk�H��$�   L�D$xH�<
I�4 �   �Hc�$�   Hk�HcL$$Hk�H�T$hH�|$HH��$  H�<
H��$  H�4�   󤋄$�   9D$(��   HcD$(H�L$X��$�   9���   �D$(��H�H�L$X���������D$0�D$(��H�H�L$X������$�   ��$�   ��$�   ��$�    t ��$�   t-��$�   t;��$�   tI�]HcD$0Hk�H�L$8�T$$��FHcD$0Hk�H�L$8�T$$�T�.HcD$0Hk�H�L$8�T$$�T�HcD$0Hk�H�L$8�T$$�T�D$(���D$(������D$$���D$$�D$p���D$p��$�   9D$(�������$�   9D$pt1L��� A�)  H��� H�Ϡ �*�  H�Ӡ �)  �	*����$�   9D$pt
�T  �O  �s  HcD$ Hk�HcL$ Hk�H�T$8H�|$8�L9LtǄ$�      �Ǆ$�       ��$�   ��$�   H�|$x �I  HcD$ Hk�H�L$8HcHk��L$$Hc�Hk�H��$�   H�|$xH��$�   H�<
H��$�   H�4�   �HcD$ Hk�H�L$8HcDHk��L$$��Hc�Hk�H��$�   H�|$xH��$   H�<
H��$   H�4�   �HcD$ Hk�H�L$8HcDHk��L$$��Hc�Hk�H��$�   H�|$xH��$P  H�<
H��$P  H�4�   󤃼$�    tQHcD$ Hk�H�L$8HcDHk��L$$��Hc�Hk�H��$�   H�|$xH��$0  H�<
H��$0  H�4�   �HcD$ Hk�H�L$8HcHk�HcL$$Hk�H�T$hH�|$HH��$p  H�<
H��$p  H�4�   �HcD$ Hk�H�L$8�T$$��D$$���D$$HcD$ Hk�H�L$8HcDHk�HcL$$Hk�H�T$hH�|$HH��$�   H�<
H��$�   H�4�   �HcD$ Hk�H�L$8�T$$�T�D$$���D$$HcD$ Hk�H�L$8HcDHk�HcL$$Hk�H�T$hH�|$HH��$  H�<
H��$  H�4�   �HcD$ Hk�H�L$8�T$$�T�D$$���D$$��$�    tkHcD$ Hk�H�L$8HcDHk�HcL$$Hk�H�T$hH�|$HH��$  H�<
H��$  H�4�   �HcD$ Hk�H�L$8�T$$�T�D$$���D$$�$HcD$ Hk�HcL$ Hk�H�T$8H�|$8�D�D
�q���H�L$X�ی��H�L$x�ь���  H��$�  �  =  ��  H��$�  ��  H��$�   H��$�  �  ��$�   �D$     �
�D$ ���D$ ��$�   9D$ }dHcD$ H��$�   �<� u��HcD$ H��$�   �|� tHcD$ H��$�   ���L$$�A�D$$�HcD$ H��$�   ���L$$�DA��D$$�HcD$DHk�H�> H�IH��$(  L�[� �Y  ��H��$(  ��P  H�D$HH�|$H u3���  D�D$DH�T$HH�L$h��  Hc�$�   H��H��= H�IH��$8  L� � �^  ��H��$8  ��P  H��$�   H��$�    u3��^  D��$�   H��$�   H��$�   �  �D$$�+���D���T$$H��$�  ������uH�L$H�	���H��$�   �����3��  H��$�  �X  H�D$hH��$�  �  H��$�   �D$,    �D$`    �D$     �
�D$ ���D$ ��$�   9D$ �  HcD$ H��$�   �<� u���D$P    �
�D$P���D$P�D$P��HcL$ H��$�   ;���   �D$,��;D$$}�D$`�L$P�D;D$D|H��� �t  �#���   �D$P�L$`ȋ�H�Hk�HcL$,Hk�H�T$hH�|$HH��$H  H�<
H��$H  H�4�   �D$,���D$,�D$`�L$P�DH�Hk�HcL$,Hk�H�T$hH�|$HH��$X  H�<
H��$X  H�4�   �D$,���D$,����HcD$ H��$�   �|� ��   �D$,��;D$$}�D$P�L$`ȋ�;D$D|H�2� �}  ��"���   �D$P�L$`ȋ�H�Hk�HcL$,Hk�H�T$hH�|$HH��$h  H�<
H��$h  H�4�   �D$,���D$,HcD$`Hk�HcL$,Hk�H�T$hH�|$HH��$x  H�<
H��$x  H�4�   �D$,���D$,HcD$ H��$�   ���L$`ȋ��D$`������D$     �
�D$ ���D$ �D$$�+���9D$ }+HcD$ H��$�   �D�    HcD$ H��$�   ��   �H��$�   �$���H�L$H�����   � H�L$H�	���H�L$x�����H�L$X�����3�H�Ĉ  _^����������L�L$ �T$�T$H�L$H��(H��9 H���   L�L$H�T$@�T$8H�L$0��  H��(������������L�L$ L�D$�T$H�L$H��(H��9 H���   L�L$HL�D$@�T$8H�L$0��   H��(��������������D�L$ L�D$�T$H�L$H��HH�J9 H���   H��$�   H�L$0H�L$xH�L$(H�L$pH�L$ D�L$hL�D$`�T$XH�L$P��(  H��H�������������D�L$ L�D$�T$H�L$H��XH��8 H���   H��$�   H�L$H��$�   �D$@H��$�   H�L$8H��$�   H�L$0H��$�   H�L$(H��$�   H�L$ D�L$xL�D$p�T$hH�L$`��0  H��X��������������D�D$H�T$H�L$H��(H�>8 H���   D�D$@H�T$8H�L$0��@  H��(���������������������̉T$H�L$H��(H��7 H���   �T$8H�L$0���  H��(�������������������\$ �T$H�T$H�L$H��XH��7 H���   ��$�   �L$@H��$�   H�L$8��$�   �L$0H��$�   H�L$(H��$�   H�L$ �\$x�T$pH�T$hH�L$`���  H��X�����������H�L$H�D$H�g� H�H�D$H�@    H�D$����������H�L$H��(H�D$0H�3� H�H��6 H���   H�L$0H�I�PH��(����������D�L$ L�D$�T$H�L$H��8H��6 H���   H�L$@H�I�PH�|$P u�   �NH��6 H���   L�L$`D�D$XH�T$P�L$H�H�L$@H�AH�D$@H�x t
�D$    ��D$     �D$ H��8��������������H�L$H��(H�D$0H�x u3��H�6 H���   H�L$0H�I�P H��(���������D�L$ D�D$�T$H�L$H��HH�D$0H�D$ L�L$4D�D$`�T$XH�L$P��  �D$h9D$4u�D$0���D$h9D$0u�D$4������H��H������������D�L$ L�D$H�T$H�L$H��HH�Y5 H���   H��$�   H�L$0H�L$xH�L$(�L$p�L$ D�L$hL�D$`H�T$XH�L$P���  H��H�������������L�L$ L�D$H�T$H�L$H��8H��4 H���   H�L$`H�L$ L�L$XL�D$PH�T$HH�L$@��  H��8�������������������\$ �T$�T$H�L$H��(WҋT$8H�L$0�V����T$H�L$@�  (ЋT$8H�L$0�$���H��(�����������������\$ �T$�T$H�L$H��   H�L$H�ra��L��D��$�   H�T$0H��$�   ��`����$�   ��$�   �D$@�  �D$ ��$�   ��$�   �D$8�m  �D$(��$�   ��$�   �D$0�J  �L$ (��L$((�(�H�L$`�`��L����$�   H��$�   �`��H�Ĉ   �������������L�L$ L�D$H�T$H�L$H��8H�93 H���   �L$`�L$ L�L$XL�D$PH�T$HH�L$@��`  H��8��������������������H�L$H�D$����������������������H�L$�����������H��(H��2 H���   ���  H��(��������������������H�L$H��(H��2 H���   H�L$0���  H��(����������L�L$ D�D$H�T$H�L$H��hH�I2 H���   H��$�   H�L$X��$�   �L$PH��$�   H�L$HH��$�   H�L$@��$�   �L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ L��$�   D��$�   H�T$xH�L$p���  H��h��������������������L�L$ D�D$H�T$H�L$H��hH��1 H���   H��$�   H�L$X��$�   �L$PH��$�   H�L$HH��$�   H�L$@��$�   �L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ L��$�   D��$�   H�T$xH�L$p���  H��h��������������������H�L$H��(H��0 H���   H�L$0��X  H��(����������H�T$H�L$H��(H��0 H���   H�T$8H�L$0���  H��(����������������H�L$H��(H�h0 H���   H�L$0���  H��(����������L�D$H�T$H�L$H��(H�.0 H���   L�D$0H�T$8H�L$@���  H��(������D�D$H�T$H�L$H��(HcD$@Hk�L��H�T$0H�L$8�7 H��(��������������D�D$H�T$H�L$H��(HcD$@H��L��H�T$0H�L$8�b7 H��(��������������L�L$ L�D$H�T$H�L$H��XH�T$xH�L$x��  ��t`H�� �7 L��� H��� H���S  H�D$@�   @�   ��   L�x� A�}  H�L$@H�ы���  �0/ ��t��fH�D$hH�L$pH��H�D$8H�T$pH�L$`�  H��H�D$ L�L$8L�D$hH�T$`H�L$0��	  H�D$pH�D$ L�L$8L�D$hH�T$`H�L$0�  H��X�����������L�D$H�T$H�L$H��(H�|$@~L�L$8L�D$@H�T$8H�L$0�����H��(�������̉T$�L$�D$�L$ȋ������������̉T$H�L$H��(H�L$0�	����D$8����t
H�L$0�j[��H�D$0H��(�����������L�D$H�T$H�L$H��8H�L$P�5 H;D$@vH�D$PH�D$ �
H�D$HH�D$ H�D$ H��8�������������H�T$H�L$H��(H��- H���   H�T$8H�L$0���  H��(�����������������T$�L$�D$�D$f/D$v�D$��D$f/D$v�D$��D$������������L�L$ L�D$H�T$H�L$H��8H�|$` ~DH�D$PH   H�D$ L�L$ L�D$PH�T$HH�L$@�  L�L$XL�D$ H�T$HH�L$@�  �%H�D$XH9D$PtL�L$XL�D$PH�T$HH�L$@�g  H��8���L�L$ L�D$H�T$H�L$H��xH��* H3�H�D$`H��$�   }��  H��$�   H�D$0H�D$0H�H+�H��H��H�D$83�����  H�|$8~H�D$8H��H�D$8�   H�D$0H��H�D$0H��$�   H�L$8H�D��H�D$PH��$�   H�L$0H��H�D$HA�   H�T$PH�L$X�s3 A�   H�T$HH�L$P�^3 A�   H�T$XH�L$H�I3 H�|$0�  H�D$8H�D$(H��$�   H�L$(H�D��H�D$ H�D$(H�H;D$0��   H�D$ H�D$@H�D$(H�H�D$(H��$�   H�L$(H�D��H�D$ H�D$0H9D$(}5H�D$ H��H��H�L$ �h  ��tH�D$(H��H�D$(H�D$ H��H�D$ H�T$ H�L$@�:  ��tAA�   H�T$@H�L$X�q2 A�   H�T$ H�L$@�\2 A�   H�T$XH�L$ �G2 ���#����R���H�L$`H3��3 H��x��������H�T$H�L$H��(H�C* H���   H�T$8H�L$0��`  H��(����������������H�L$H�D$�@���H�L$H��(H��) H���   H�L$0�PXH��(�������������L�L$ D�D$�T$H�L$H��8H��) H���   H�L$`H�L$ L�L$XD�D$P�T$HH�L$@H�I�PH��8���H�L$H��8H�D$@�x ~�   Hk� H�L$@HH����  �D$ ��D$ �����D$ H��8�������������H�L$H��(H�() H��  H�L$0���   H��(����������H�L$H��(H��( H��  H�L$0�PPH��(�������������H�L$H��(��  H�L$0�8  H��(����H�L$H��(E3���  H�L$0�  H��(ÉT$H�L$H��(H��( H���   �T$8H�L$0H�I�P(H��(�H�L$H��(��  H�L$0��   H��(����H�L$H��(E3���  H�L$0��   H��(�H�L$H��(E3���  H�L$0��   H��(�H�L$H��(�(  H�L$0�h   H��(����H�L$H��(E3��(  H�L$0�   H��(�D�D$�T$H�L$H��(H��' H���   D�D$@�T$8H�L$0��(  H��(�������̉T$H�L$H��(H�t' H���   �T$8H�L$0��8  H��(��D�D$�T$H�L$H��(H�?' H���   D�D$@�T$8H�L$0���  H��(��������D�D$�T$H�L$H��(H��& H���   D�D$@�T$8H�L$0��0  H��(��������H�L$H��(H��& H��  H�L$0�PH��(������������̉T$H�L$H��(HcD$8H�L$0H�	H��H���
   H��(������H�L$H�D$� %���3ҹ   ��������H�T$H�L$H��(H�C& H��  H�T$8H�L$0���   H��(����������������L�L$ L�D$H�T$H�L$H��XH�Q$ H3�H�D$@H�D$pH�L$xH+�H��H��H�� ~0H�D$pH�L$xH+�H��H��L��L�D$pH�T$hH�L$`�4�����   H�D$pH��H�D$0H�D$0H�D$ H�D$ H��H�D$(�H�D$ H��H�D$ H�D$(H��H�D$(H�D$pH9D$ tTH�T$(H�L$ ��  ��tAA�   H�T$ H�L$8��, A�   H�T$(H�L$ ��, A�   H�T$8H�L$(��, �H�D$0H��H�D$0H�D$xH9D$0�L���H�L$@H3�� . H��X������������L�L$ L�D$H�T$H�L$H��XH�D$pH�L$xH+�H��H��H�� ��   H��$�    uL�L$xL�D$pH�T$hH�L$`�V�����   H��$�   H��H��$�   H�D$xH��H�D$8H�L$pH�T$xH+�H��H��H��H�H+�H��H�L$pH��H�L$8H�L$ L��L�D$pH�T$hH�L$`�  H�D$@H�D$@H�D$ L�L$xL�D$pH�T$hH�L$`�o  H�D$0H��$�   H�D$ L�L$xL�D$0H�T$hH�L$`�����H�D$0H�D$x�����H��XÉT$H�L$H��(H��# H���   �T$8H�L$0��x  H��(�̉T$H�L$H��(HcD$8H�L$0H�	H��H���
   H��(������H�L$H��H�D$ � %   ���u	�$   ��$    �$H�����������������̉T$H�L$H��(H��" H���   �T$8H�L$0�PXH��(�����D�D$�T$�L$�D$9D$}�D$��D$9D$~�D$��D$���������������H�T$H�L$H��H�D$ H�L$(�	9}	�$   ��$    �$H�������������H�T$H�L$H��H�$    �H�D$(H��H�D$(H�|$(tH�$H��H�$��H�$H����������������L�L$ L�D$H�T$H�L$H��(H�T$HH�L$@�I�����t?H�T$PH�L$H�6�����t	H�D$H�`�H�T$PH�L$@������tH�D$P�DH�D$@�=�6H�T$PH�L$@�������t	H�D$@�!�H�T$PH�L$H�������tH�D$P�H�D$HH��(�������L�D$�T$H�L$H��(H�/! H��  L�D$@�T$8H�L$0�P H��(�����������D�D$H�T$H�L$H��(H��  H���   D�D$@H�T$8H�L$0�PPH��(���������H�T$H�L$H��(H��  H��  H�T$8H�L$0���   H��(����������������L�L$ L�D$H�T$H�L$H��(�H�D$@H��H�D$@H�D$HH9D$@tL�D$@H�T$8H�L$0�   ��H��(��L�D$H�T$H�L$H��HH�v H3�H�D$0H�D$`H��H��H�L$`�x�����txA�   H�T$`H�L$(�' H�D$(H�D$ H�D$`H��A�   H��H�L$`�' H�D$`H��H�D$`H�D$`H��H��H�L$ ������u�A�   H�T$ H�L$`�L' H�L$0H3��( H��H�����������L�L$ L�D$H�T$H�L$H��8H�� H3�H�D$(H�D$PH��H�D$P3�����   H�D$PH��H�D$PH�T$`H�L$P������t��H�D$XH��H�D$XH�T$XH�L$`�`�����t��H�D$XH9D$PrH�D$P�rA�   H�T$PH�L$ �& A�   H�T$XH�L$P�m& A�   H�T$ H�L$X�X& H�D$`H9D$PuH�D$XH�D$`�H�D$`H9D$Xu
H�D$PH�D$`�*���H�L$(H3��x' H��8����L�L$ L�D$H�T$H�L$VWH��H  H��$p   u$H��$h  H��$`  �   �H��$h  �5  H��$`  L��$x  H��H�L$H�G   H��$`  �@P�D$@�|$@ t1�|$@��   �|$@��  �|$@��  �|$@��  �  H��$`  H��L��$x  H��H��$X  �l#  H��$�   H��$`  L��$x  H��H��$�  �  H�D$8    H�D$0    H��$�  �A�D$(H��$�  ��D$ H��$�   L��L��H��$  H��$p  � H�L$HH��H��   ���  H��$`  H��L��$x  H��H��$h  �"  H�D$xH��$`  L��$x  H��H��$8  ��  H�L$hH�L$0H��$�  �A�D$(H��$�  ��D$ H�L$xL��L��H��$  H��$p  � H�L$HH��H��   �|$h �V  �f W�W�H��$h  �GI��H��$�   H��$`  L��$x  H��H��$  �K  L��H��$�  H��$p  �#(  H��$�   H��$`  H��H��$`  L��H��$H  �7   L��$x  H��H��$�  ��  L��H��$�  H��$p  ��'  H��$�   L��H��H��$�  �l  H��H��$x  ��  H��$�   L��H��H��$�   �a   H��$`  L��$x  H��H��$(  �q  H��$�   H��$`  L��$x  H��H��$8  �I  L��H��$�   H��$p  �!'  L��$�   H��H��$�  �I  L��H��$�  H��$p  �%  H��$�   L��H��H��$�  �  H��H��$�  �  H��$�   H��H��   �H��$`  L��$x  H��H��$�  �  H�D$8    H�D$0    H��$�  �A�D$(H��$�  ��D$ L��$�   L��H��$�   H��$p  � H�L$HH��H��   ���  H��$�  �@f.nv zt1L��$�  H��$�   H��$p  �$  H�L$HH��H��   ��oL�D$HH��$   H��$p  �o%  �XH��$�  �PH��$�  �H��$P  �xF��L��H��$�  H��$p  �<$  H�L$HH��H��   ��  H��$`  H��L��$x  H��H��$�  ��  H��$�   H��$`  H��0L��$x  H��H��$�  �%  H�D$0    H��$�  �A�D$(H��$�  ��D$ H��$�   L��L��H��$  H��$p  �� H�L$HH��H��   �H��$`  H��0L��H�T$HH��$@  �Q  H��H��$p  ��  L��H��$`  �HHH��$�  �  H��$`  H��0L��H��H��$�  �  H�L$HH��H��   ���  H��$`  H��0L��$x  H��H��$   �  A�   H��H��$p  �� H��$`  �HH�Y�(��D$`�D$`f.,t zu��w �D$`H��$`  H��0L��$x  H��H��$0  �  L��H��$`  H��$p  �~#  L��H��$�  H��$�  �&  H�L$HH��H��   �W��D$XH�L$H�Q!  �L$`�  �D$pH�T$HH��$�  �^  L���L$pH��$�  �X  H�L$HH��H��   ��D$p�^D$`�5  ��  fWw �YD$`�D$XH��$`  H��0L��$x  H��H��$   �  L��H��$P  H��$p  �"  L��H�T$HH��$�  �  L��H��$�  H��$p  �#!  H�L$HH��H��   �H��$x  H��$�  �  L��H�T$HH��$h  �7  H��$h  H��H  _^����������������������L�L$ L�D$H�T$H�L$������������L�L$ D�D$H�T$H�L$H��  H�D$@������$   t
�   ��  H��$�   �B��H��$  H� H��$  H��$  ���   �D$(�|$( u
�   �  H��$(  H��$  ��  �D$0H��$0  ��  H�D$8�/   H�L$H�+X  �   H�L$`�X  L�D$8H��$  H��$(  �   �D$     �
�D$ ���D$ �|$ �  �|$  uE3�H�T$`H��$(  �   �E3�H�T$HH��$(  �    �D$$    �
�D$$���D$$�D$(9D$$��   �D$09D$$u
�D$,   ��D$,    �D$ 9D$,t��H��$�   �)  �H��$  H� L��$�   D�D$$H��$  H��$  ���   ��$�   �uH��$�   �s	  �h���E3�A�   H��$�   H��$(  ��  �H��$�   �B	  �7���������   H��  ������������L�L$ L�D$H�T$H�L$�   �������D�L$ L�D$H�T$H�L$H��  H�D$(�����   ��$H  �+  ��t
������%  H��$�   H��$(  �8  �D$$�����D$     �
�D$ ���D$ H��$   H� H��$(  H��$   ���   9D$ ��   H�L$0��  �H��$   H� L�L$0D�D$ H��$(  H��$   ���   ��$�   �uH�L$0�  �|���L��$�   H�T$0H��$�   �  D��$@  D��$8  H��H��$0  ��  ��t)�D$ �D$$�   ��$H  �  ��uH�L$0�  �H�L$0�  �����D$$H��  �����������������L�L$ L�D$H�T$H�L$VWH��  H�D$H����H��$�  �=  H�D$@H��$P  H��$�  �  H�L$@L��H��H��$�   ��  H�L$p�  �3�H��$�  �!  H�D$8H�D$8H� L�L$pD��$�  H��$�  H�L$8���   H��$�  H�D$ L��$�   L��$   H��$�   H�L$p����H�L$PH��H��   �H��$�  H� H�L$pH�L$ L�L$PD��$�  H��$�  H��$�  ��   �D$0   H�L$p�I  �D$0H�ĸ  _^������������L�D$H�T$H�L$3����������������L�L$ L�D$H�T$H�L$3�����������L�L$ L�D$H�T$H�L$������������L�D$H�T$H�L$3����������������L�L$ L�D$H�T$H�L$�   �������L�D$H�T$H�L$������������������\$ L�D$H�T$H�L$3����������L�L$ L�D$H�T$H�L$������������H�T$H�L$3���������������������L�L$ D�D$H�T$H�L$������������L�L$ D�D$H�T$H�L$������������L�L$ D�D$H�T$�L$H��x  H��$�  ��  ��t"E3�H��$�  ��$�  �nl����u3���   E3��@  H�L$0����H�D$(    H��$�  H�D$ D��$�  D��$�  H��$�  H�L$0�   H��  H��$�  ��$�  ����tH��  H��$�  ��$�  �� ��tH��  H��$�  ��$�  %�   ��tH��  H��$�  ��$�  ����tH�d  H��$�  �D$ @  L�L$0L��$�  ��$�  �   �^H  H��x  �������D�L$ D�D$H�T$H�L$H��8H�D$hH�D$(�D$X�D$ L�L$`L�D$H�T$PH�L$@�����H�D$@H�L$`H��@  H�D$@H�i  H��H  H�D$@H�b  H��P  H�D$@H�[  H���  H�D$@H�T  H��X  H�D$@H�M  H���  H�D$@H�R  H���  H�D$@H�3  H���  H�D$@H�8  H���  H��8�H�L$VWH��xH��$�   H���:��H��$�   H��H����9��H��$�   H��0H����9��W�H�L$ 耎��H�D$ H��$�   H��   �W�H�L$8�\���H��$�   H�L$8H�xH��   �W�H�L$P�4���H��$�   H�L$PH�x0H��   �H��$�   ��h �@HH��$�   �@P    H��$�   H��x_^������̉T$H�L$H��(H�D$0�T$8H���r  H�D$0H���T$8H���]  H�D$0H��0�T$8H���H  H�D$0H��H�T$8H���3  H�D$0H��(����������H�L$VWH��   H��$�   H���8��H��$�   H��H���8��H��$�   H��0H���8��H��$�   H��HH���n8��W�W�W�H�L$ �G8��H��$�   H��   �W�W���T H�L$8�8��H��$�   H�yH��   �W���T W�H�L$P��7��H��$�   H�y0H��   ���T W�W�H�L$h��7��H��$�   H�yHH��   �H��$�   H�Ĉ   _^�����̉T$H�L$H�D$��H�L$�����������H�T$H�L$VWH��   3�H�L$0�1���H��$�   H��$�   �@8�YAXH��$�   H��$�   �HP�YI@�\�H��$�   �H�Y�(�H��$�   H��$�   �HP�YI(H��$�   H��$�   �P �YQX�\�H��$�   �P0�Y�(��X�H��$�   H��$�   �H �YI@H��$�   H��$�   �P8�YQ(�\�H��$�   �PH�Y�(��X��D$ �D$ f.�e zuH��$�   ����H��$�   �  ��R �^D$ �D$ H��$�   H��$�   �@�YAXH��$�   H��$�   �HP�YI�\�H��$�   �H0�Y�(�H��$�   H��$�   �H�YI8H��$�   H��$�   �P�YQ@�\�H��$�   �PH�Y�(��X�H��$�   H��$�   �HP�YI@H��$�   H��$�   �P8�YQX�\�H��$�   ��Y�(��X��YD$ �D$0H��$�   H��$�   �@�YA(H��$�   H��$�   �H �YI�\�H��$�   �HH�Y�(�H��$�   H��$�   �H �YIXH��$�   H��$�   �PP�YQ(�\�H��$�   ��Y�(��X�H��$�   H��$�   �HP�YIH��$�   H��$�   �P�YQX�\�H��$�   �P�Y�(��X��YD$ �D$8H��$�   H��$�   �@8�YA(H��$�   H��$�   �H �YI@�\�H��$�   ��Y�(�H��$�   H��$�   �H@�YIH��$�   H��$�   �P8�YQ�\�H��$�   �P�Y�(��X�H��$�   H��$�   �H�YI H��$�   H��$�   �P�YQ(�\�H��$�   �P0�Y�(��X��YD$ �D$@H��$�   H��$�   �@8�YAXH��$�   H��$�   �HP�YI@�\��YD$ �D$HH��$�   H��$�   �@P�YA(H��$�   H��$�   �H �YIX�\��YD$ �D$PH��$�   H��$�   �@ �YA@H��$�   H��$�   �H8�YI(�\��YD$ �D$XH��$�   H��$�   �@@�YAHH��$�   H��$�   �HX�YI0�\��YD$ �D$`H��$�   H��$�   �@X�YAH��$�   H��$�   �H(�YIH�\��YD$ �D$hH��$�   H��$�   �@(�YA0H��$�   H��$�   �H@�YI�\��YD$ �D$pH��$�   H��$�   �@0�YAPH��$�   H��$�   �HH�YI8�\��YD$ �D$xH��$�   H��$�   �@H�YA H��$�   H��$�   �H�YIP�\��YD$ ��$�   H��$�   H��$�   �@�YA8H��$�   H��$�   �H0�YI �\��YD$ ��$�   H�D$0H��$�   H��`   �H��$�   H�Ę   _^��������H�T$H�L$H��8H�D$HH�L$H� �YH�D$HH�L$H�H�YI�X�H�D$HH�L$H�H�YI�X���  �D$ �D$ f.�_ zuW�H�L$@����H�D$@�g��L �^D$ �D$ H�D$H�@�YD$ H�D$H�H�YL$ H�D$H��YT$ �T$((�(��D$((�H�L$@��/��H�D$@H��8����L�D$H�T$H�L$VWH��   3�H�L$ �l���H��$�   H��$�   �@�YH��$�   ��X�(�H��$�   H��$�   �H0�YI�X�H��$�   H��$�   �HH�YI�X��D$ H��$�   H��$�   �@ �YH��$�   �H�X�(�H��$�   H��$�   �H8�YI�X�H��$�   H��$�   �HP�YI�X��D$(H��$�   H��$�   �@(�YH��$�   �H�X�(�H��$�   H��$�   �H@�YI�X�H��$�   H��$�   �HX�YI�X��D$0H��$�   H��$�   �@�YAH��$�   H��$�   �H0�YI �X�H��$�   H��$�   �HH�YI(�X��D$8H��$�   H��$�   �@ �YAH��$�   H��$�   �H8�YI �X�H��$�   H��$�   �HP�YI(�X��D$@H��$�   H��$�   �@(�YAH��$�   H��$�   �H@�YI �X�H��$�   H��$�   �HX�YI(�X��D$HH��$�   H��$�   �@�YA0H��$�   H��$�   �H0�YI8�X�H��$�   H��$�   �HH�YI@�X��D$PH��$�   H��$�   �@ �YA0H��$�   H��$�   �H8�YI8�X�H��$�   H��$�   �HP�YI@�X��D$XH��$�   H��$�   �@(�YA0H��$�   H��$�   �H@�YI8�X�H��$�   H��$�   �HX�YI@�X��D$`H��$�   H��$�   �@�YAHH��$�   H��$�   �H0�YIP�X�H��$�   H��$�   �HH�YIX�X��D$hH��$�   H��$�   �@ �YAHH��$�   H��$�   �H8�YIP�X�H��$�   H��$�   �HP�YIX�X��D$pH��$�   H��$�   �@(�YAHH��$�   H��$�   �H@�YIP�X�H��$�   H��$�   �HX�YIX�X��D$xH�D$ H��$�   H��`   �H��$�   H�Ĉ   _^������������L�D$H�T$H�L$H��8H�D$PH�L$H�@(�YH�D$P�H�X�(�H�D$PH�L$H�H@�YI�X�H�D$PH�L$H�HX�YI�X�H�D$PH�L$H�H �Y	H�D$P�P�X�(�H�D$PH�L$H�P8�YQ�X�H�D$PH�L$H�PP�YQ�X�H�D$PH�L$H�P�YH�D$P��X�(�H�D$PH�L$H�X0�YY�X�H�D$PH�L$H�XH�YY�X��T$ (�(��D$ (�H�L$@�)��H�D$@H��8����������L�D$�L$H�L$H��8H�D$P�@�YD$HH�D$P�H�YL$HH�D$P��YT$H�T$ (�(��D$ (�H�L$@�2)��H�D$@H��8�����L�D$H�T$H�L$H��8H�D$HH�L$P�@�\AH�D$HH�L$P�H�\IH�D$HH�L$P��\�T$ (�(��D$ (�H�L$@�(��H�D$@H��8�����������L�D$H�T$H�L$H��8H�D$HH�L$P�@�XAH�D$HH�L$P�H�XIH�D$HH�L$P��X�T$ (�(��D$ (�H�L$@�8(��H�D$@H��8����������̉T$�L$�D$�L$#ȋ�������������L�D$H�T$H�L$H��8H�D$HH�L$P� �YAH�D$HH�L$P�H�Y	�\�H�D$HH�L$P�H�Y	H�D$HH�L$P��YQ�\�H�D$HH�L$P�P�YQH�D$HH�L$P�X�YY�\��T$ (�(��D$ (�H�L$@�R'��H�D$@H��8�����L�D$H�T$H�L$H��8H�D$PH�L$H�@(�YH�D$PH�L$H�H@�YI�X�H�D$PH�L$H�HX�YI�X�H�D$PH�L$H�H �Y	H�D$PH�L$H�P8�YQ�X�H�D$PH�L$H�PP�YQ�X�H�D$PH�L$H�P�YH�D$PH�L$H�X0�YY�X�H�D$PH�L$H�XH�YY�X��T$ (�(��D$ (�H�L$@�I&��H�D$@H��8����H����   ���H����   ���H����   ���H����   ���H����   ���H����   ���H����   ���H����   ���H����   ���H����   ���H����   ���H����   ���H����   ����������������D$H��(�D$0f/0B r��X �'���X f/D$0r
��X ��D$0�U H��(�H�L$H��8H�L$@荃����t
�D$    ��D$     �D$ H��8����������������D$H��(�D$0� H��(�������D�L$ D�D$H�T$H�L$H��(H��� H���   D�L$HD�D$@H�T$8H�L$0��  H��(�������������L$�D$�D$f/D$v�D$��D$��������H�T$H�L$H��(H�� H���   H�T$8H�L$0��@  H��(����������������H�L$H��(H��� H���   H�L$0�PxH��(�������������H�T$H�L$VWH��   H��� H���   H�T$ H��$�   �PXH��$�   H��`   �H��$�   H�Ĉ   _^������������H�L$H��(H�H� H���   H�L$0�PHH��(������������̉T$H�L$H��(H�� H���   �T$8H�L$0�PpH��(�����H�T$H�L$VWH��   H��� H���   H�T$ H��$�   �PxH��$�   H��`   �H��$�   H�Ĉ   _^������������H�L$H��(H�D$0H�L$0� �YH�D$0H�L$0�H�YI�X�H�D$0H�L$0�H�YI�X��0  H��(������������D�L$ D�D$H�T$H�L$H��(H�� H���   D�L$HD�D$@H�T$8H�L$0�P(H��(���������������L�D$H�T$H�L$VWH��HH��� H���   L�D$pH�T$`H�L$ �P`H�|$hH��   �H�D$hH��H_^�L�D$H�T$H�L$H��(H�~� H���   L�D$@H�T$8H�L$0���   H��(������D�D$H�T$H�L$H��(H�>� H���   D�D$@H�T$8H�L$0�P0H��(����������D$H��(�D$0�W�  H��(�������L�D$H�T$H�L$VWH��HH��� H���   L�D$pH�T$`H�L$ �PpH�|$hH��   �H�D$hH��H_^�L�D$H�T$H�L$VWH��HH��� H���   L�D$pH�T$`H�L$ �PXH�|$hH��   �H�D$hH��H_^�H�T$H�L$H��H�D$(H�L$ �	9t3��  H�D$(�x uOH�D$(�8 uEH�D$(�x u:H�D$ �x uH�D$ �8 uH�D$ �x u	�$   ��$    �$�   �XH�D$ �x uMH�D$ �8 uCH�D$ �x u8H�D$(�x uH�D$(�8 uH�D$(�x u
�D$   ��D$    �D$�]H�D$(�x t!H�D$ �x tH�D$(H�L$ �I9Ht3��1H�D$(�x t!H�D$ �x tH�D$(H�L$ �I9Ht3���   H����������H�T$H�L$H��8H�T$HH�L$@������u
�D$    ��D$     �D$ H��8���������������������H�L$H��8��   ��  H�D$ H�|$  tH�D$ H���    u�H�L$@H�D$ ���   H�D$@H��8����������������������H�T$H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u�H�L$@H�D$ ���   H�T$HH�L$@��  H�D$@H��8�����������������̉T$H�L$H��H��   �)  H�D$ H�|$  tH�D$ H���    u�+H�L$PH�D$ ���   �T$XH�L$(�  H��H�L$P��  H�D$PH��H�������H�T$H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u�H�L$@H�D$ ���   H�T$HH�L$@�{  H�D$@H��8������������������L�D$H�T$H�L$H��8��   �C  H�D$ H�|$  tH�D$ H���    u�.H�L$@H�D$ ���   H�T$HH�L$@�  H�T$PH�L$@�W  H�D$@H��8��������������L�L$ L�D$H�T$H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u�=H�L$@H�D$ ���   H�T$HH�L$@�   H�T$PH�L$@��   H�T$XH�L$@��   H�D$@H��8����������H�L$H��8��   �=  H�D$ H�|$  tH�D$ H���    u�H�L$@H�D$ ���   H��8�����������H�T$H�L$H��8��   ��  H�D$ H�|$  tH�D$ H���    u�H�T$HH�L$@H�D$ ���   H��8�����������������H�T$H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u�H�T$HH�L$@H�D$ ���   H��8�����������������H�L$H��8��   �-  H�D$ H�|$  tH�D$ H���    u�H�L$@H�D$ ���   H��8����������̉T$H�L$H��8��   ��  H�D$ H�|$  tH�D$ H���    u	H�V� ��T$HH�L$@H�D$ ���   H��8������������H�T$H�L$H��8��   �x  H�D$ H�|$  tH�D$ H���    uH�D$@�H�T$@H�L$HH�D$ ���   H�D$@H��8�������H�T$H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u3��H�T$@H�L$HH�D$ ���   H��8���������������H�T$H�L$H��8��   �  H�D$(H�|$( tH�D$(H���    u�   �/H�T$@H�L$HH�D$(���   ��u
�D$    ��D$     �D$ H��8������������������D�D$H�T$H�L$H��hH�D$@�����D$     ��   �"  H�D$(H�|$( tH�D$(H���    u$H��� H�L$x�%�����D$ ���D$ H�D$x�UD��$�   H�T$pH�L$HH�D$(���   H�D$0H�D$0H�D$8H�T$8H�L$x������D$ ���D$ H�L$H�B���H�D$xH��h���������H�T$H�L$H��8�x  �h  H�D$ H�|$  tH�D$ H��x   u3��H�T$HH�L$@H�D$ ��x  H��8���������������H�T$H�L$H��8�x  �  H�D$ H�|$  tH�D$ H���   u3��H�T$HH�L$@H�D$ ���  H��8���������������H�L$H��8�D$     �
�D$ ���D$ �T$ H�L$@�����8 t��D$ H��8����������������������L�D$H�T$H�L$H��8�D$     �
�D$ ���D$ �T$ H�L$@�K����8 t9�T$ H�L$H�8���H�D$(�T$ H�L$@�%���H�L$(H��H��������t��H�|$P tH�D$P�L$ ��|$  ~�T$ H�L$@������8 u
�D$$   ��D$$    �D$$H��8����������������������H�T$H�L$H��H��  �  H�D$ H�|$  tH�D$ H���   uH�D$P�)L�D$XH�T$PH�L$(H�D$ ���  H�L$(�����H�D$PH��H��������L�D$H�T$H�L$H��hH�D$@�����D$     ��  �  H�D$(H�|$( tH�D$(H���   u"H�T$xH�L$p�'�����D$ ���D$ H�D$p�UL��$�   H�T$xH�L$HH�D$(���  H�D$0H�D$0H�D$8H�T$8H�L$p������D$ ���D$ H�L$H�$���H�D$pH��h�����������H�L$H�D$����������������������H��8�   �2  H�D$ H�|$  tH�D$ H�x u3��H�D$ �PH��8���������H�L$H��8H�D$@H�8 u�>�   ��  H�D$ H�|$  tH�D$ H�x u�H�L$@H�D$ �PH�D$@H�     H��8��������D�D$H�T$H�L$H��8H�|$H u3��>�    �w  H�D$ H�|$  tH�D$ H�x  u3��D�D$PH�T$HH�L$@H�D$ �P H��8��������������̉T$H�L$H��8�(   �  H�D$ H�|$  tH�D$ H�x( u3���T$HH�L$@H�D$ �P(H��8�������H�T$H�L$H��8�0   ��  H�D$ H�|$  tH�D$ H�x0 u3��H�T$HH�L$@H�D$ �P0H��8���������������������H�L$H��8�8   �m  H�D$ H�|$  tH�D$ H�x8 u3��H�L$@H�D$ �P8H��8���������������H�L$H��8�@   �  H�D$ H�|$  tH�D$ H�x@ u3��H�L$@H�D$ �P@H��8���������������L�L$ L�D$H�T$H�L$H��8�H   �  H�D$ H�|$  tH�D$ H�xH u3��L�L$XL�D$PH�T$HH�L$@H�D$ �PHH��8�����������������L�D$H�T$H�L$H��8�P   �S  H�D$ H�|$  tH�D$ H�xP u3��L�D$PH�T$HH�L$@H�D$ �PPH��8�����������L�L$ L�D$H�T$H�L$H��8�H   ��
  H�D$ H�|$  tH�D$ H�xX u3��L�L$XL�D$PH�T$HH�L$@H�D$ �PXH��8�����������������H�L$H��8�`   �
  H�D$ H�|$  tH�D$ H�x` u3��H�L$@H�D$ �P`H��8���������������L�L$ L�D$H�T$H�L$H��H�h   �.
  H�D$0H�|$0 tH�D$0H�xh u3��&H�D$pH�D$ L�L$hL�D$`H�T$XH�L$PH�D$0�PhH��H�������H�T$H�L$H��8�p   ��	  H�D$ H�|$  tH�D$ H�xp u�H�T$HH�L$@H�D$ �PpH��8�������H�T$H�L$H��8�P  �x	  H�D$ H�|$  u3��H�T$HH�L$@H�D$ ��P  H��8��������������H�T$H�L$H��8�X  �(	  H�D$ H�|$  u3��H�T$HH�L$@H�D$ ��X  H��8��������������H�T$H�L$H��8�`  ��  H�D$ H�|$  u3��H�T$HH�L$@H�D$ ��`  H��8��������������L�L$ L�D$H�T$H�L$H��8�h  �~  H�D$ H�|$  u�L�L$XL�D$PH�T$HH�L$@H�D$ ��h  H��8������������H�L$H��8��   �-  H�D$ H�|$  tH�D$ H���    u3��H�L$@H�D$ ���   H��8���������H�T$H�L$H��8��   ��  H�D$ H�|$  u�H�T$HH�L$@H�D$ ���   H��8����������������H�T$H�L$H��8��   �  H�D$ H�|$  u3��H�T$HH�L$@H�D$ ���   H��8��������������L�D$�T$H�L$H��8��   �4  H�D$ H�|$  u3��L�D$P�T$HH�L$@H�D$ ���   H��8����������������������L�L$ L�D$H�T$H�L$H��8�H  ��  H�D$ H�|$  u3��L�L$XL�D$PH�T$HH�L$@H�D$ ��H  H��8����������L�L$ L�D$H�T$H�L$H��H�@  �n  H�D$0H�|$0 u3��3H�D$xH�D$(H�D$pH�D$ L�L$hL�D$`H�T$XH�L$PH�D$0��@  H��H����������������������H�L$H��8��   ��  H�D$ H�|$  u3��H�L$@H�D$ ���   H��8��������H�T$H�L$H��8��   �  H�D$ H�|$  u�H�T$HH�L$@H�D$ ���   H��8����������������L�D$H�T$H�L$H��xH�D$@�����D$     ��   �R  H�D$(H�|$( tH�D$(H���    u23�H�L$H�Z  H��H��$�   �J�����D$ ���D$ H��$�   �^L��$�   H�T$XH��$�   H�D$(���   H�D$0H�D$0H�D$8H�T$8H��$�   �����D$ ���D$ H�L$X�^���H��$�   H��x������������������L�L$ L�D$H�T$H�L$H��8��  �n  H�D$ H�|$  tH�D$ H���   u3��L�L$XL�D$PH�T$HH�L$@H�D$ ���  H��8�����������H�T$H�L$H��8�  �  H�D$ H�|$  tH�D$ H��   u3��H�T$HH�L$@H�D$ ��  H��8���������������H�T$H�L$H��8�  �  H�D$ H�|$  tH�D$ H��   u3��H�T$HH�L$@H�D$ ��  H��8���������������H�T$H�L$H��8�  �H  H�D$ H�|$  tH�D$ H��   u3��H�T$HH�L$@H�D$ ��  H��8���������������H�L$H��8�   ��  H�D$ H�|$  tH�D$ H��    u3��H�L$@H�D$ ��   H��8���������L�L$ L�D$H�T$H�L$H��8�(  �  H�D$ H�|$  tH�D$ H��(   u3��L�L$XL�D$PH�T$HH�L$@H�D$ ��(  H��8�����������H�T$H�L$H��8�0  �(  H�D$ H�|$  tH�D$ H��0   u�H�T$HH�L$@H�D$ ��0  H��8�����������������L�L$ D�D$H�T$H�L$H��8�8  �  H�D$ H�|$  tH�D$ H��8   u3��L�L$XD�D$PH�T$HH�L$@H�D$ ��8  H��8�����������H�L$H��8��  �]  H�D$(H�|$( tH�D$(H���   u3��H�L$@H�D$(���  �D$ �D$ H��8�����������������L�D$H�T$�L$H��8�   ��   H�D$ H�|$  tH�D$ H�x u3��L�D$PH�T$H�L$@H�D$ �PH��8�������������H�T$H�L$H��hH�D$@�����D$     �h  �   H�D$(H�|$( uH�L$p�����D$ ���D$ H�D$p�MH�T$xH�L$HH�D$(��p  H�D$0H�D$0H�D$8H�T$8H�L$p�
���D$ ���D$ H�L$H�@��H�D$pH��h�����������̉L$H��(L��� �T$0�D ���  H��(��������������̉T$H�L$H�D$�L$�H�D$�@    H�D$�@    H�D$���������������D�L$ D�D$H�T$�L$H��X�   ��  H�D$@H�|$@ tH�D$@H�x u������<��$�   �D$0��$�   �D$(��$�   �D$ D�L$xD�D$pH�T$h�L$`H�D$@�PH��X���������������D�L$ D�D$H�T$�L$H��   H�D$`�����   �c  H�D$HH�|$H tH�D$HH�x u�D$D����H��$�   �%D���D$D�{H�D$hH�D$PH��$�   H�L$P�C��H�D$X��$�   �D$0��$�   �D$(��$�   �D$ D��$�   D��$�   H�T$X��$�   H�D$H�P�D$@H��$�   �C���D$@H�Ę   �������������H�T$�L$H��8�   �   H�D$ H�|$  tH�D$ H�x u3��H�T$H�L$@H�D$ �PH��8������̉L$H��8�    �>   H�D$ H�|$  tH�D$ H�x  u3���L$@H�D$ �P H��8����������������̉L$H��(L�� �T$0��f �3�  H��(���������������H�L$H�D$H��� H��� � ������D�D$H�T$H�L$H��8H��� H��  H�L$@���   H�D$ H�|$  u3��D�D$PH�T$HH�L$ �o  H��8�����������D�D$H�T$H�L$H��8H�^� H��  H�L$@���   H�D$ H�|$  u3��D�D$PH�T$HH�L$ �O  H��8�����������H�T$H�L$H��(H�D$0H�L$8H�H��� H�@ E3�E3�3�H�L$0H�	�P H�L$0H�AH�D$0H��(���������������������H�L$H��(H��� H�@ E3�E3�3�H�L$0H�	�P H�L$0H�AH��(������������L�D$H�T$H�L$H��(H�D$0H�x u3��7H�N� H�@ H�L$0L�IL�D$@H�T$8H�L$0H�	�P H�L$0H�A�   H��(��D�D$H�T$H�L$H��(H��� H���   D�D$@H�T$8H�L$0�PH��(���������D�D$H�T$H�L$H��(H��� H���   D�D$@H�T$8H�L$0�PpH��(���������L�L$ L�D$H�T$�L$H��h�D$p�D$ �|$ t7�|$ �#  �|$ �  �|$ t�|$ ��   �  �   �}  �U� ���M� �=F� ��   H�L$x����=�6  }
������G  H��$�    u
������2  L�I5 A�m   H��� �(   �,��H�D$(H�|$( tH�L$(��=��H�D$0�	H�D$0    H�D$0H�D$@H�D$@H��� H�=��  tH��$�   H��� ��D���   �   H��$�   �L$x�� ����u
������   �   �   �l ����W� �ȉO� �=H�  u\������6��H�=,�  t=H�#� H�D$HH�D$HH�D$8H�|$8 t�   H�L$8�=6��H�D$P�	H�D$P    H���     �   ������H��h������������������L�D$�T$H�L$H���D$(�$�<$t�H�D$ H��� H�D$0H�� �   H����������������H�L$H��(H�H� H�@ E3������H�L$0�P(H�D$0H��(������������������̉T$H�L$H��(H�� H�@ E3��T$8H�L$0�P(H�D$0H��(����������������H�T$H�L$H��(H��� H�@ L�D$8�����H�L$0�P(H�D$0H��(������������H�L$H��(H�L$0�  H��(���������H�T$H�L$H��(E3�E3�H�T$0H�L$8�-  H�D$0H��(��������������������H�T$H�L$H��(H�#� H�@ H�T$8H�L$0�PH��(����������������������H�T$H�L$H��8H��� H�@ H�T$HH�L$@�P��u
�D$    ��D$     �D$ H��8������������L�D$�T$H�L$H��(A�#  L�D$@�T$8H�L$0�e  H��(�����������������L�D$�T$H�L$H��(A�F  L�D$@�T$8H�L$0�%  H��(����������������̉T$H�L$H��8�T$HH�L$@��  H�D$ H�L$ �V  H��8������������������D�D$�T$H�L$H��8�T$HH�L$@�  H�D$ �T$PH�L$ �=  H��8��������̉T$H�L$H��8H��� H�@ �T$HH�L$@���  H�D$ H�|$  u3��
H�L$ ��\��H��8����������H�T$H�L$H��(H�C� H�@ H�T$8H�L$0���  H��(���L�L$ D�D$H�T$H�L$H��(H�	� H�@ L�L$HD�D$@H�T$8H�L$0��   H��(���������������H�L$H��(H��� H�@ H�L$0�P8H��(����������������H�L$H��(H��� H��  H�L$0���   H��(���������̉T$H�L$H��(H�d� H��  �T$8H�L$0���   H��(�̉T$H�L$H��(H�4� H�@ �T$8H�L$0���   H��(�����D�L$ L�D$�T$H�L$H��(H��� H�@ D�L$HL�D$@�T$8H�L$0���   H��(�H�L$H��(H�D$0H��(H���6/  H��(������������������H�T$H�L$H��(H��� H�@pH�T$8H�L$0���   H��(�������������������H��(H�]� H�@p�PxH��(����������H�L$H��(H�8� H�@pH�L$0H�	���   H�D$0H�     H��(��������������L�L$ L�D$H�T$H�L$H��HH��� H�@p��$�   �L$0�L$x�L$(�L$p�L$ L�L$hL�D$`H�T$XH�L$P�PH��H�������L�L$ L�D$H�T$H�L$H��8H��� H�@p�L$h�L$(�L$`�L$ L�L$XL�D$PH�T$HH�L$@�PH��8������������������H��(H�=� H�@p�H��(�����������H�L$H��(H�� H�@pH�L$0H�	�PH�D$0H�     H��(�����������������D�L$ L�D$H�T$H�L$H��(H��� H�@pD�L$HL�D$@H�T$8H�L$0�P H��(������������������D�D$H�T$H�L$H��(H�~� H�@pD�D$@H�T$8H�L$0�P0H��(������������H�L$H��(H�H� H�@pH�L$0�P8H��(����������������H�T$H�L$H��(H�� H�@pH�T$8H�L$0�P@H��(����������������������D�L$ L�D$H�T$H�L$H��8H��� H�@p�L$h�L$(�L$`�L$ D�L$XL�D$PH�T$HH�L$@�PHH��8������������������L�D$H�T$H�L$H��(H�n� H�@pL�D$@H�T$8H�L$0�PPH��(������������L�L$ L�D$H�T$H�L$H��(H�)� H�@pL�L$HL�D$@H�T$8H�L$0�PXH��(������������������D�L$ L�D$H�T$H�L$H��(H��� H�@pD�L$HL�D$@H�T$8H�L$0�P(H��(������������������L�D$H�T$H�L$H��(H��� H�@pL�D$@H�T$8H�L$0�P`H��(������������L�L$ L�D$H�T$H�L$H��(H�I� H�@pL�L$HL�D$@H�T$8H�L$0�PhH��(������������������H�T$H�L$H��(H�� H�@pH�T$8H�L$0�PpH��(����������������������H�T$�L$H��XH�D$hH��xH�L$hH��`H�T$hH��HL�D$hI��0L�L$hI��L�L$@L�T$hL��� M�[H�D$0H�L$(H�T$ M��H�D$@L��I�ҋL$`A��p  H��X���������������������H��(H�=� H�@��x  H��(�������H��(H�� H�@���  H��(������̉L$H��(H��� H�@�L$0�PXH��(������������������L�L$ D�D$�T$�L$H��HH��� H�@H��$�   H�L$0H�L$xH�L$(H�L$pH�L$ L�L$hD�D$`�T$X�L$P��@  H��H������������������H�L$H��XH�D$(�����D$     H�L$0�:����H�<� H�@H�L$0�PpH�T$0H�L$`�I����D$ ���D$ H�L$0����H�D$`H��X�����������H��(H��� H�@�PxH��(���������̉T$H�L$H��(H��� H�@�T$8H�L$0���   H��(���������������������H��(H��� H�@���   H��(�������H��(H�m� H�@���   H��(�������L�D$H�T$H�L$H��(H�>� H�@L�D$@H�T$8H�L$0���   H��(��������̉T$H�L$H��(H�� H�@�T$8H�L$0���   H��(���������������������H�L$H��(H��� H�@H�L$0��x  H��(�������������H�L$H��(H��� H�@H�L$0��X  H��(�������������L�L$ L�D$�T$�L$H��8H�[� H�@�L$`�L$(H�L$XH�L$ L�L$PD�D$H�T$@��6  ��h  H��8����������������H�L$H��(H�� H�@H�L$0�PH��(����������������H�L$H��xH�D$0����E3�H��& H�L$P�&���H�D$ H�D$ H�D$(L��$�   H�T$(H�L$8�H���H�L$P����H��� H�@H�L$8�P�H�L$8�����H��x�������L�D$H�T$H�L$H��(H�N� H�@L�D$@H�T$8H�L$0��   H��(���������H�L$H��(H�� H�@H�L$0��p  H��(�������������H�L$H��hH�D$8�����D$     H��� H�@H�L$@��  H�D$(H�D$(H�D$0H�T$0H�L$p������D$ ���D$ H�L$@����H�D$pH��h��������������������H�L$H��hH�D$8�����D$     H�W� H�@H�L$@��  H�D$(H�D$(H�D$0H�T$0H�L$p�R����D$ ���D$ H�L$@����H�D$pH��h��������������������D�L$ D�D$H�T$H�L$H��(H��� H�@D�L$HD�D$@H�T$8H�L$0���  H��(��������������̉T$H�L$H��(H��� H�@�T$8H�L$0���  H��(��������������������̉T$�L$H��(H�U� H�@�T$8�L$0��   H��(������̉T$�L$H��(H�%� H�@�T$8�L$0��  H��(������̉L$H��(H��� H�@�L$0��  H��(��������������̉L$H��(H��� H�@�L$0���   H��(���������������H�L$H��(H��� H�@H�L$0���   H��(�������������H�L$H��(H�h� H�@H�L$0���   H��(�������������H��(H�=� H�@���   H��(������̉L$H��(H�� H�@�L$0��(  H��(���������������H��(H��� H�@���   H��(�������H��(H��� H�@���   H��(������̉L$H��(H��� H�@�L$0���   H��(���������������H�L$H��(H�x� H�@H�L$0���   H��(�������������D�D$�T$�L$H��(H�@� H�@D�D$@�T$8�L$0���   H��(������������̉L$H��(H�	� H�@�L$0���  H��(���������������D�L$ D�D$�T$�L$H��(H�˿ H�@D�L$HD�D$@�T$8�L$0��  H��(�������������������H�T$�L$H��(H��� H�@H�T$8�L$0���   H��(���������������������H�T$�L$H��(H�D� H�@H�T$8�L$0���  H��(��������������������̉T$H�L$H��hH�D$(�����D$     H�L$0�)���H�� H�@H�T$0�L$x���   H�T$0H�L$p�*���D$ ���D$ H�L$0�y*��H�D$pH��h����������������H�T$�L$H��(H��� H�@H�T$8�L$0��   H��(���������������������L�L$ L�D$H�T$H�L$H��(H�9� H�@L�L$HL�D$@H�T$8H�L$0���  H��(���������������H�T$H�L$H��(H�� H�@H�T$8H�L$0���  H��(�������������������L�D$H�T$H�L$H��(H��� H�@L�D$@H�T$8H�L$0��  H��(���������H��(H�}� H�@��  H��(�������H�L$H��XH�D$(�����D$     H�L$0������H�<� H�@H�L$0��  H�T$0H�L$`�F����D$ ���D$ H�L$0�q���H�D$`H��X��������H��(H�� H�@���  H��(�������H�L$H��(H�ȼ H�@H�L$0��  H��(������������̉T$H�L$VWH��HH��� H�@�T$hH�L$ ��`  H�|$`H��   �H�D$`H��H_^�������������H�T$�L$H��(H�D� H�@H�T$8�L$0��H  H��(���������������������D�L$ �T$�L$�L$H��(H��� H�@D�L$H�T$@�L$8�L$0��  H��(�������������D�D$H�T$�L$H��(H��� H�@D�D$@H�T$8�L$0���  H��(�����������D�D$H�T$�L$H��(H�o� H�@D�D$@H�T$8�L$0���  H��(�����������D�D$H�T$�L$H��(H�/� H�@D�D$@H�T$8�L$0���  H��(�����������D�D$H�T$�L$H��(H�� H�@D�D$@H�T$8�L$0���  H��(����������̉L$H��(H��� H�@�L$0��   H��(���������������D�D$H�T$�L$H��(H�� H�@D�D$@H�T$8�L$0��  H��(����������̉T$H�L$H��(H�D� H�@�T$8H�L$0���  H��(���������������������H��(H�� H�@���  H��(�������L�L$ L�D$H�T$�L$H��(H�ڹ H�@L�L$HL�D$@H�T$8�L$0���  H��(�����������������D�L$ D�D$H�T$H�L$H��8H��� H�@H�L$`H�L$ D�L$XD�D$PH�T$HH�L$@���  H��8��������������������̉L$H��(H�9� H�@�L$0���  H��(���������������H�L$H��(H�� H�@H�L$0���  H��(�������������H�L$H��(H�ظ H�@H�L$0���  H��(������������̉T$H�L$H��hH�D$8�����D$     H��� H�@�T$xH�L$@��(  H�D$(H�D$(H�D$0H�T$0H�L$p�����D$ ���D$ H�L$@�����H�D$pH��h�����������̉T$H�L$H��hH�D$8�����D$     H�� H�@�T$xH�L$@��0  H�D$(H�D$(H�D$0H�T$0H�L$p�
����D$ ���D$ H�L$@�@���H�D$pH��h������������H�L$H��(H��� H�@H�L$0��8  H��(�������������H�L$H��(H�x� H�@H�L$0��@  H��(�������������H�L$H��8H�H� H�@L�L$(L�D$$H�T$ H�L$@���  ��u3���D$ H��8������������������H�L$H��8H��� H�@L�L$(L�D$ H�T$$H�L$@���  ��u3���D$ H��8������������������H�L$H��8H��� H�@L�L$(L�D$ H�T$$H�L$@���  ��u3��H�D$(H��8�����������������L�D$�T$�L$H��(H�P� H�@L�D$@�T$8�L$0���  H��(������������̉T$�L$H��(H�� H�@�T$8�L$0���  H��(������̉T$�L$H��(H�� H�@�T$8�L$0���  H��(������̉L$H��(H��� H�@�L$0���  H��(��������������̉L$H��(H��� H�@�L$0���  H��(���������������H�L$H��(H�X� H�@H�L$0���  H��(�������������H�T$�L$H��(H�$� H�@H�T$8�L$0��   H��(��������������������̉L$H��(H�� H�@�L$0���  H��(��������������̉T$H�L$H��xH�D$8�����D$     H��� H�@��$�   H�L$@���  H�D$(H�D$(H�D$0H��$�   H�L$0�D!���D$ ���D$ H�L$@� ��H��$�   H��x�������������������H�L$H��(H�(� H�@H�L$0���  H��(������������̉L$H��(H��� H�@�L$0���  H��(���������������H��(H�ͳ H�@���  H��(������̉L$H��(H��� H�@�L$0��p  H��(���������������H�L$H�T$L�D$L�L$ H��H  H��� H3�H��$0  H��$X  H�D$ L�L$ L��$P  �   H�L$0��  H�+� H�@H�T$0H�� ��h  H�D$     H��$0  H3��$�  H��H  �������������H�L$H��83�H�L$@蛩  H�D$ H�|$  tH�L$ �4���H�L$ � ��H��8����������������������D�L$ D�D$H�T$H�L$H��hH�L$x�Η��H�o� H�I`H�L$P��$�   �T$H��$�   �T$@��$�   �T$8��$�   �T$0��$�   �T$(��$�   �T$ D��$�   D��$�   H��H�L$pH�D$P��p  H��h���������������������D�L$ D�D$H�T$H�L$H��hH�L$x�n  H��� H�I`H�L$P��$�   �T$H��$�   �T$@��$�   �T$8��$�   �T$0��$�   �T$(��$�   �T$ D��$�   D��$�   H��H�L$pH�D$P��p  H��h���������������������D�L$ D�D$H�T$H�L$H��XH�� H�@`��$�   �L$H��$�   �L$@��$�   �L$8��$�   �L$0��$�   �L$(��$�   �L$ D�L$xD�D$pH�T$hH�L$`��p  H��X�������������H�L$H��(H��� H�@`H�L$0��h  H��(�������������D�D$�T$H�L$H��(H�_� H�@`D�D$@�T$8H�L$0��`  H��(�����������L�L$ L�D$H�T$H�L$H��8H�� H�@`H�L$`H�L$ L�L$XL�D$PH�T$HH�L$@��x  H��8���������������������H�L$H��(H�ȯ H�@`H�L$0��X  H��(�������������L�L$ L�D$H�T$H�L$H��8H��� H�@`H�L$`H�L$ L�L$XL�D$PH�T$HH�L$@���  H��8���������������������H��(H�=� H�@`��H  H��(�������H�L$H��(H�� H�@`H�L$0H�	��P  H�D$0H�     H��(��������������D�L$ L�D$�T$H�L$H��XH�D$8�����D$     H��� H�@D�L$xL�D$p�T$hH�L$@���  H�D$(H�D$(H�D$0H�T$0H�L$`�F����D$ ���D$ H�L$@�1���H�D$`H��X��������H�L$H��xH�D$8�����D$     �LGOgH�L$P����H�D$(H�D$(H�D$0E3�L�D$0�icMCH�L$@�!����H�L$P�f���H�L$@�\��H��u,H��$�   �����D$ ���D$ H�L$@蕍��H��$�   �7H�L$@�!��H��H��$�   ������D$ ���D$ H�L$@�\���H��$�   H��x����������������H�L$H��(H�h� H�@H�L$0��`  H��(�������������D�L$ D�D$�T$�L$H��HH�+� H�@H��$�   H�L$8H��$�   H�L$0�L$x�L$(H�L$pH�L$ D�L$hD�D$`�T$X�L$P��h  H��H�������D�L$ D�D$�T$�L$H��XH��� H�@��$�   �L$@H��$�   H�L$8H��$�   H�L$0��$�   �L$(��$�   �L$ D�L$xD�D$p�T$h�L$`���  H��X��������D�L$ D�D$H�T$H�L$H��xH�D$H�����D$0    H�(� H�@H�D$(    ��$�   �L$ D��$�   D��$�   H��$�   H�L$P���  H�D$8H�D$8H�D$@H�T$@H��$�   ������D$0���D$0H�L$P�*���H��$�   H��x�������������������D�L$ D�D$H�T$H�L$H��hH�D$H�����D$0    H�h� H�@H��$�   H�L$ D��$�   D��$�   H�T$xH�L$P���  H�D$8H�D$8H�D$@H�T$@H�L$p�����D$0���D$0H�L$P�̊��H�D$pH��h������������������̉T$�L$H��XH�D$ �����������u�d���H�L$8�����D�D$`���H�L$8�w���D�D$h���H�L$8�c���E3�L�D$8�icMCH�L$(����H�L$(�7����H�L$8�����H��X�������̉T$H�L$H��xH�D$8�����D$     �]�����u&H��$�   ������D$ ���D$ H��$�   �   �!��H�L$P������D��$�   �!��H�L$P����E3�L�D$P�icMCH�L$@�����H�D$(H�D$(H�D$0H�L$0����H��H��$�   ������D$ ���D$ H�L$@�W����H�L$P�����H��$�   H��x���������������̉T$H�L$H��xH�D$8�����D$     �m�����u&H��$�   �*�����D$ ���D$ H��$�   �   ����H�L$P������D��$�   ����H�L$P�����E3�L�D$P�icMCH�L$@�����H�D$(H�D$(H�D$0H�L$0����H��H��$�   ������D$ ���D$ H�L$@�g����H�L$P�����H��$�   H��x���������������̉L$H��xH�D$8����������u3��t�#��H�L$P�3����D��$�   �#��H�L$P����E3�L�D$P�icMCH�L$@�4���H�D$(H�D$(H�D$0H�L$0軍���D$ H�L$@轇���H�L$P�R����D$ H��x���������̉L$H��xH�D$8�����������u3��t�s��H�L$P�����D��$�   �s��H�L$P�f���E3�L�D$P�icMCH�L$@����H�D$(H�D$(H�D$0H�L$0�����D$ H�L$@�����H�L$P�����D$ H��x����������D�L$ L�D$�T$�L$H��8H�� H�@H�L$hH�L$(�L$`�L$ D�L$XL�D$P�T$H�L$@��x  H��8�����������������D�L$ D�D$H�T$H�L$H��8H��� H�@H�L$hH�L$(�L$`�L$ D�L$XD�D$PH�T$HH�L$@���  H��8�������������L�D$H�T$H�L$H��(H�^� H�@L�D$@H�T$8H�L$0���  H��(���������H�L$H��(H�D$0H�8 tH�� H�@H�L$0H�	���  H�D$0H�     H��(�������������������H�L$H��(H�إ H�@H�L$0���  H��(�������������H�L$H��(H��� H�@H�L$0���  H��(�������������D�D$H�T$H�L$H��(H�n� H�@D�D$@H�T$8H�L$0���  H��(���������D�D$H�T$H�L$H��(H�.� H�@D�D$@H�T$8H�L$0���  H��(���������D�D$H�T$H�L$H��(H�� H�@D�D$@H�T$8H�L$0���  H��(���������D�D$H�T$H�L$H��(H��� H�@D�D$@H�T$8H�L$0���  H��(���������H��(H�}� H�@���  H��(�������L�L$ L�D$H�T$H�L$H��HH�I� H�@��$�   �L$0H�L$xH�L$(H�L$pH�L$ L�L$hL�D$`H�T$XH�L$P���  H��H����������������H�T$H�L$H��(H�� H�@H�T$8H�L$0���  H��(�������������������L�L$ D�D$H�T$H�L$H��(H��� H�@L�L$HD�D$@H�T$8H�L$0���  H��(���������������H��(H�]� H�@���  H��(�������L�D$�T$H�L$H��(H�/� H�@L�D$@�T$8H�L$0���  H��(�����������H��(H��� H�@���  H��(�������H��(H�ݢ H�@��  H��(������̉T$H�L$H��hH�D$8�����D$     H��� H�@�T$xH�L$@��  H�D$(H�D$(H�D$0H�T$0H�L$p�����D$ ���D$ H�L$@�����H�D$pH��h������������H�L$H��(H�8� H�@H�L$0��  H��(������������̉L$H��(H�	� H�@�L$0��   H��(��������������̉T$H�L$H��(H�ԡ H�@�T$8H�L$0��(  H��(���������������������H�L$H��(H��� H�@H�L$0��0  H��(�������������D�D$H�T$�L$H��(H�_� H�@D�D$@H�T$8�L$0��8  H��(�����������D�D$H�T$H�L$H��(H�� H�@D�D$@H�T$8H�L$0��@  H��(���������D�D$�T$�L$H��(H�� H�@D�D$@�T$8�L$0���  H��(�������������L�D$H�T$H�L$H��(H��� H�@L�D$@H�T$8H�L$0��`  H��(���������H�L$H��(H�h� H�@H�L$0��H  H��(������������̉T$H�L$H��(H�4� H�@�T$8H�L$0��H  H��(���������������������H�L$H��(H��� H�@H�L$0��P  H��(�������������H�L$H��(H�ȟ H�@H�L$0��X  H��(�������������H��(H��� H�@��`  H��(�������H��(H�}� H�@��x  H��(�������D�L$ D�D$�T$�L$H��HH�K� H�@H��$�   H�L$8H��$�   H�L$0�L$x�L$(�L$p�L$ D�L$hD�D$`�T$X�L$P��  H��H���������L�D$H�T$�L$H��(H�ߞ H�@L�D$@H�T$8�L$0���  H��(�����������H�L$H��(H��� H�@H�L$0���  H��(�������������H�L$H��(H�x� H��  H�L$0��  H��(����������H�L$H�D$H�@��L�L$ L�D$�T$H�L$H��8�|$H 3��kHcD$HL�L$XL�D$PH��H�L$@� �D$ �|$  |�D$H��9D$ |3�|$  }H�� �H  �B����D$H��H�H�L$@� �D$H�ȉD$ �D$ H��8���������������H�L$H��XH�D$`� �i  �D$8H�D$`�@�T  �D$0�.� f/D$8w�� f/D$0v#H�D$`W�� H�D$`�-� �@��  �� f/D$8��   �� f/D$0��   �,D$8�D$$�,D$0�D$ �|$  u H�D$`W�� H�D$`��� �@�f�D$$��|$ �D$(�D$ �D$$�D$(�D$ �|$( u��*D$$H�D$`��^�(�H�D$`� �*D$$H�D$`�H�^�(�H�D$`�@�-  �L$0�D$8�L  �� �^�(��D$@�'� f/D$@vV�D$8�YD$@�D$8�D$0�YD$@�D$0H�D$`� �YD$@H�D$`� H�D$`�@�YD$@H�D$`�@��� f/D$0v ��� �D$0H�D$`��� �@�L$0�D$8��  �D$H�D$0�D$8�D$H�D$0�D$Hf/�  s�H�D$`� �^D$8H�D$`� H�D$`�@�^D$8H�D$`�@H��X�������������L$H�L$H��(�D$8f/�  v��  �D$8��  f/D$8v�{  �D$8�D$8�Y�� �X?  �*$��H�D$0� H�D$0��� �@H�L$0�����H�D$0H��(�������������T$�L$H�L$H��8�D$Hf/� r
�D$$   ��D$$    �D$Pf/�� r
�D$    ��D$     �D$ 9D$$u
�D$(   ��D$(    �D$(�D$,�D$H��  �Xp� �[#��H�D$@� �D$P�  �XO� �:#��H�D$@�@H�D$@��� f/@v#H��� �   ����H�D$@��� �@�|$, uH�D$@� fW� H�D$@� H�L$@����H�D$@H��8����������������������L$H�L$H��(H�D$0�D$8�@H�D$0�� f/@v#H�6� �,   �l���H�D$0��� �@H��(�����������������������L$H�L$H��8��� f/D$HvH�� �5   ������� �D$HH�D$@� �YD$H��!���D$ H�D$@�@��!���L$ �^�(���!��H�D$@� �D$H�!��H�D$@�@H�L$@����H��8������������D$H��(�D$0�m�  H��(��������L$�D$�D$f/D$v�D$��D$���������L$�D$H��(�L$8�D$0��  H��(�����������H�L$H��(H�D$0H� H�L$0�PH��(�������������������H�L$H��(H�D$0H� H�L$0�PH��(�������������������H�L$H��(H�D$0H��� H�H�D$0�@    H�� H���   L�'  L�D$0H�����H�T����H�L$0H�AH�D$0H��(����������������H�L$H��(H�D$0H�k� H�H�D$0�x uH��� H���   H�L$0H�I�PH��(���������������D�D$�T$H�L$H��(H�D$0H�x u3��&H�_� H���   E3�D�D$@�T$8H�L$0H�I�PH��(�������������������̉T$H�L$H��(H�D$0H�x tH�� H���   �T$8H�L$0H�I�PH��(��������������������̉T$H�L$H��(H�D$0H�x tH��� H���   �T$8H�L$0H�I�P H��(���������������������H�L$H�D$H�     H�D$�@    H�D$��������������H�L$H��(H�D$0H�8 u�AH�;� H���   H�L$0H�	���   H�� H���   H�L$0H�	�PxH�D$0H�     H��(���������������������L�L$ D�D$H�T$H�L$H��HH�D$PH�8 t1H��� H���   H�L$PH�	�PxH�D$PH�     H�D$P�@    H�D$P�L$`�HH��� H���   H��  H�L$(H�L$hH�L$ L�����L������T$`H�L$X�PpH�L$PH��D$0    �
�D$0���D$0�D$`9D$0��   HcD$0H�L$hH���x uBHcD$0H�L$hH���@   HcD$0H�L$hH��H�� H���   H�L$8H�HH�D$8�PH�Ó H���   �T$0H�L$PH�	���   HcL$0H�T$hH��H�A�[���H�D$PH�8 t
�D$4   ��D$4    �D$4H��H����������������������L�L$ D�D$H�T$H�L$H��(H�L$8�  L�L$HD�D$@H��H�L$0�7���H��(������������������̉T$H�L$H��8H�D$(    �D$     �
�D$ ���D$ H�D$@�@9D$ }yH�ɒ H���   �T$ H�L$@H�	���   H�D$(H�|$( t'H��� H���   E3�D�D$H�   H�L$(�P��u H�u� H���   H�L$@H�	���   3��
�o����   H��8����������������������H�L$H��(H�(� H���   H�L$0H�	���   H��(�������H�L$H��(H��� H���   H�L$0H�	���   H��(�������H�L$H��(H�ȑ H���   H�L$0H�	���   H��(�������H��(H��� H���   ���   H��(��������������������H�L$H��(H�h� H���   H�L$0���   H��(����������H��(H�=� H���   ��  H��(��������������������H�L$H��(H�� H���   H�L$0��  H��(����������H�L$H��(H�D$0H� H�L$0�PH��(��̉T$H�L$H��(H�L$0������D$8����t
H�L$0�
���H�D$0H��(�����������H�L$H�D$H�@��H�L$3����������H�L$H��(H�X� H���   H�L$0��@  H��(����������L�D$H�T$H�L$H��(H�� H���   L�D$@H�T$8H�L$0��H  H��(����������������������H�T$H�L$H��8H�ӏ H���   H�L$@��@  H�D$ H�|$  u#H��� H���   E3�H�T$HH�L$@��H  �H�L$ �?2  H��H�L$H�"i��H��8��������������H�L$H��(H�X� H���   H�L$0��P  H��(����������L�D$H�T$H�L$H��(H�� H���   L�D$@H�T$8H�L$0��X  H��(����������������������H��(H�ݎ H���   �H��(��������H�L$H��(H��� H���   H�L$0H�	�P H�D$0H�     H��(��������������H��(H�}� H���   ���  H��(��������������������H�L$H��(H�H� H���   H�L$0H�	�P H�D$0H�     H��(��������������D�D$H�T$H�L$H��hH�D$8�����D$     H�� H���   D��$�   H�T$pH�L$@�PH�D$(H�D$(H�D$0H�T$0H�L$x�ۻ���D$ ���D$ H�L$@����H�D$xH��h�������������L�D$�T$H�L$H��(H�o� H���   L�D$@�T$8H�L$0�P H��(����������̉T$H�L$H��(H�4� H���   �T$8H�L$0���  H��(������������������H�L$H��(H��� H���   H�L$0�P(H��(�������������H�L$H��(H�Ȍ H���   H�L$0�P0H��(�������������H�L$H��(H��� H���   H�L$0�P8H��(�������������L�L$ L�D$H�T$H�L$H��(H�Y� H���   L�L$HL�D$@H�T$8H�L$0�P@H��(���������������H�T$H�L$H��(H�� H���   H�T$8H�L$0��h  H��(����������������D�L$ L�D$H�T$H�L$H��(H�ɋ H���   D�L$HL�D$@H�T$8H�L$0�PHH��(���������������L�L$ L�D$H�T$H�L$H��8H�y� H���   �L$`�L$ L�L$XL�D$PH�T$HH�L$@�PPH��8�������H�L$H��(H�8� H���   H�L$0�PXH��(�������������H�L$H��(H�� H���   H�L$0�P`H��(�������������H�L$H��(H�؊ H���   H�L$0�PhH��(�������������H�L$H��(H��� H���   3�H�L$0�PpH��(�����������L�D$H�T$H�L$H��(H�n� H���   L�D$@H�T$8H�L$0��0  H��(����������������������D�D$H�T$H�L$H��(H�� H���   D�D$@H�T$8H�L$0��   H��(����������������������D�D$H�T$H�L$H��(H�Ή H���   D�D$@H�T$8H�L$0���  H��(����������������������D�L$ D�D$H�T$H�L$H��8H�y� H���   �L$`�L$ D�L$XD�D$PH�T$HH�L$@���  H��8��������������������H�T$H�L$H��(H�#� H���   H�T$8H�L$0��(  H��(����������������H�T$H�L$H��(H�� H���   H�T$8H�L$0��P  H��(����������������H�T$H�L$H��(H��� H���   H�T$8H�L$0���  H��(����������������D�D$H�T$H�L$H��(H�^� H���   D�D$@H�T$8H�L$0��  H��(����������������������D�D$H�T$H�L$H��(H�� H���   D�D$@H�T$8H�L$0��`  H��(����������������������D�D$H�T$H�L$H��(H��� H���   D�D$@H�T$8H�L$0��h  H��(����������������������H�T$H�L$H��(H�s� H���   H�T$8H�L$0�PxH��(�������������������D�D$H�T$H�L$H��(H�.� H���   D�D$@H�T$8H�L$0���  H��(����������������������H�L$H��(H�� H���   H�L$0�PH��(�������������D�D$�T$H�L$H��(H��� H���   D�D$@�T$8H�L$0���   H��(��������H�T$H�L$H��(H�s� H���   E3�H�T$8H�L$0���   H��(�������������H�T$H�L$H��(H�3� H���   A�   H�T$8H�L$0���   H��(����������H�T$H�L$H��(H�� H���   E3�H�T$8H�L$0���   H��(�������������H�T$H�L$H��(H��� H���   A�   H�T$8H�L$0���   H��(����������H�L$H��(H�x� H���   H�L$0��8  H��(����������L�D$H�T$H�L$H��hH�D$8�����D$     H�-� H���   L��$�   H�T$pH�L$@��  H�D$(H�D$(H�D$0H�T$0H�L$x�����D$ ���D$ H�L$@�C���H�D$xH��h����������H�L$H��xH�D$0����H�L$H�t�����  H�L$8����H��H�L$X�����E3�L�D$HH�T$XH��$�   �+����u
�D$$   ��D$$    �D$$�D$ H�L$X�C����D$ ��t�D$(    H�L$H��c���D$(�H�L$H��i���D$,H�L$H��c���D$,H��x������������������H�L$H��hH�D$ �����   H�L$H�?�����  H�L$(�?���H��H�L$8�2����A�   L�D$HH�T$8H�L$p�7+���H�L$8茔���H�L$H�Qc��H��h�������������H�T$H�L$H��xH�D$0�����D$$    H�L$H������  H�L$8跩��H��H�L$X誒���E3�L�D$HH�T$XH��$�   �_*����u
�D$(   ��D$(    �D$(�D$ H�L$X�����D$ ��t,H��$�   � ����D$$���D$$H�L$H�b��H��$�   �7H�L$H�%  H��H��$�   ������D$$���D$$H�L$H�Rb��H��$�   H��x����������������������H�T$H�L$H��xH�D$0�����D$$    H�L$H������  H�L$8觨��H��H�L$X蚑���E3�L�D$HH�T$XH��$�   �O)����u
�D$(   ��D$(    �D$(�D$ H�L$X�֒���D$ ��t,H��$�   ������D$$���D$$H�L$H�{a��H��$�   �7H�L$H��#  H��H��$�   ������D$$���D$$H�L$H�Ba��H��$�   H��x����������������������H�T$H�L$H��hH�D$ ����H�T$xH�L$H�!  ���  H�L$(蚧��H��H�L$8荐���A�   L�D$HH�T$8H�L$p�(���H�L$8�����H�L$H�`��H��h��������H�T$H�L$H��hH�D$ ����H�T$xH�L$H�*!  ���  H�L$(����H��H�L$8�����A�   L�D$HH�T$8H�L$p�(���H�L$8�g����H�L$H�,`��H��h��������H�L$H��xH�D$8����H�L$P������  H�L$@褦��H��H�L$`藏���E3�L�D$PH�T$`H��$�   �L'����u
�D$$   ��D$$    �D$$�D$ H�L$`�Ӑ���D$ ��tW��D$(H�L$P�_���D$(� H�L$P�"  �D$0H�L$P�e_���D$0H��x������������L$H�L$H��hH�D$ �����L$xH�L$H�(   ���  H�L$(�ȥ��H��H�L$8軎���A�   L�D$HH�T$8H�L$p��&���H�L$8�����H�L$H��^��H��h����������������������H�L$H��xH�D$0����H�L$H� �����  H�L$8�D���H��H�L$X�7����E3�L�D$HH�T$XH��$�   ��%����u
�D$$   ��D$$    �D$$�D$ H�L$X�s����D$ ��t�D$(    H�L$H�(^���D$(�H�L$H�d���D$,H�L$H�
^���D$,H��x�����������������̉T$H�L$H��hH�D$ �����T$xH�L$H�������  H�L$(�l���H��H�L$8�_����A�   L�D$HH�T$8H�L$p�d%���H�L$8蹎���H�L$H�~]��H��h����������H�T$H�L$VWH��hH�D$(����H�L$@�M������  H�L$0����H��H�L$P������E3�L�D$@H�T$PH��$�   �$����u
�D$$   ��D$$    �D$$�D$ H�L$P�����D$ ��t"H��$�   �����H�L$@��\��H��$�   �.H�L$@�   H��$�   H��   �H�L$@�\��H��$�   H��h_^�������������H�T$H�L$H��hH�D$ ����H�T$xH�L$H�  ���  H�L$(�����H��H�L$8�����A�   L�D$HH�T$8H�L$p��#���H�L$8�G����H�L$H�\��H��h��������H�T$H�L$VWH��hH�D$(����H�L$@��������  H�L$0�}���H��H�L$P�p����E3�L�D$@H�T$PH��$�   �%#����u
�D$$   ��D$$    �D$$�D$ H�L$P謌���D$ ��t"H��$�   �����H�L$@�[[��H��$�   �.H�L$@�  H��$�   H��   �H�L$@�+[��H��$�   H��h_^�������������H�T$H�L$H��hH�D$ ����H�T$xH�L$H�J  ���  H�L$(芡��H��H�L$8�}����A�   L�D$HH�T$8H�L$p�"���H�L$8�׋���H�L$H�Z��H��h��������L�D$H�T$H�L$VWH��8H��z H���   A�   L�D$`H�T$PH�L$ ���  H�|$XH��   �H�D$XH��8_^��������L�D$H�T$H�L$VWH��8H�Lz H���   E3�L�D$`H�T$PH�L$ ���  H�|$XH��   �H�D$XH��8_^�����������H�T$H�L$VWH��hH�D$(����H�L$@�������  H�L$0�M���H��H�L$P�@����E3�L�D$@H�T$PH��$�   �� ����u
�D$$   ��D$$    �D$$�D$ H�L$P�|����D$ ��t"H��$�   �v����H�L$@�+Y��H��$�   �.H�L$@�g  H��$�   H��   �H�L$@��X��H��$�   H��h_^�������������H�T$H�L$H��hH�D$ ����H�T$xH�L$H�  ���  H�L$(�Z���H��H�L$8�M����A�   L�D$HH�T$8H�L$p�R ���H�L$8觉���H�L$H�lX��H��h��������H�T$H�L$VWH��hH�D$(����H�L$@�=������  H�L$0�ݞ��H��H�L$P�Ї���E3�L�D$@H�T$PH��$�   �����u
�D$$   ��D$$    �D$$�D$ H�L$P�����D$ ��t"H��$�   �����H�L$@�W��H��$�   �.H�L$@��  H��$�   H��   �H�L$@�W��H��$�   H��h_^�������������H�T$H�L$H��hH�D$ ����H�T$xH�L$H�  ���  H�L$(����H��H�L$8�݆���A�   L�D$HH�T$8H�L$p�����H�L$8�7����H�L$H��V��H��h��������H�L$H��xH�D$0����H�L$H��������  H�L$8�t���H��H�L$X�g����E3�L�D$HH�T$XH��$�   �����u
�D$$   ��D$$    �D$$�D$ H�L$X裇���D$ ��t�D$(    H�L$H�XV���D$(�H�L$H�8\���D$,H�L$H�:V���D$,H��x�����������������̉T$H�L$H��hH�D$ �����T$xH�L$H�������  H�L$(蜜��H��H�L$8菅���A�   L�D$HH�T$8H�L$p����H�L$8�����H�L$H�U��H��h����������H�T$H�L$VWH��hH�D$(����H�L$@�}������  H�L$0����H��H�L$P�����E3�L�D$@H�T$PH��$�   ������u
�D$$   ��D$$    �D$$�D$ H�L$P�L����D$ ��t"H��$�   �F����H�L$@��T��H��$�   �.H�L$@�7  H��$�   H��   �H�L$@��T��H��$�   H��h_^�������������H�T$H�L$H��hH�D$ ����H�T$xH�L$H��  ���  H�L$(�*���H��H�L$8�����A�   L�D$HH�T$8H�L$p�"���H�L$8�w����H�L$H�<T��H��h��������H�L$H��xH�D$0����H�L$H�������  H�L$8贚��H��H�L$X觃���E3�L�D$HH�T$XH��$�   �\����u
�D$$   ��D$$    �D$$�D$ H�L$X�����D$ ��t�D$(    H�L$H�S���D$(�H�L$H�xY���D$,H�L$H�zS���D$,H��x�����������������̉T$H�L$H��hH�D$ �����T$xH�L$H�������  H�L$(�ܙ��H��H�L$8�ς���A�   L�D$HH�T$8H�L$p�����H�L$8�)����H�L$H��R��H��h����������H�L$H��xH�D$0����H�L$H��������  H�L$8�d���H��H�L$X�W����E3�L�D$HH�T$XH��$�   �����u
�D$$   ��D$$    �D$$�D$ H�L$X蓃���D$ ��t�D$(    H�L$H�HR���D$(�H�L$H�(X���D$,H�L$H�*R���D$,H��x�����������������̉T$H�L$H��hH�D$ �����T$xH�L$H�������  H�L$(茘��H��H�L$8�������   �   �  D��L�D$HH�T$8H�L$p�x���H�L$8�͂���H�L$H�Q��H��h��������������H�L$H��8H�L$@�=����D$ �|$ t�|$ t�|$ t
�D$$    ��D$$   �D$$H��8����������H�L$H��(H�Xq H���   H�L$0���   H��(����������H�L$H��(H�(q H���   H�L$0���   H��(����������D�L$ L�D$�T$H�L$H��(H��p H���   D�L$HL�D$@�T$8H�L$0��   H��(��������������H�T$H�L$H��(H��p H���   H�T$8H�L$0��8  H��(���������������̉T$H�L$H��(H�dp H���   �T$8H�L$0���  H��(������������������H�L$H��(H�(p H���   H�L$0���   H��(����������D�L$ L�D$H�T$H�L$H��(H��o H���   D�L$HL�D$@H�T$8H�L$0���   H��(�����������̉T$H�L$H��   HǄ$�   �����/  H�D$(H�|$( u3���  H�D$8    H�D$0    H�D$     H��$�   �����H�L$P�H  �H�D$(H�D$PH��$�   H�D$`D��$�   �]  H��$�   �����E3�E3�H�T$(H��$�   �  ��u��   H�L$(�����H�D$ �
H�D$8H�D$ H�|$  ��   H�L$ ��E��H�D$8H�D$ H�D$XH�T$P��   �V�����u�   H�|$x u�   3�H�L$x�  H�D$0H�|$0 u�nH�T$ H�L$0�  H�L$x�����H�|$  tH�Un H���   H�L$ �P H�D$     �L���H�D$(H�D$@H�L$P�L����H��$�   �~���H�D$@�WH�|$( tH� n H���   H�L$(�P H�D$(    H�L$x�V���H�D$H    H�L$P�����H��$�   �%���H�D$HH�Ĩ   ���������H�L$H��(H��m H���   H�L$0���   H��(����������H�L$H��(H�hm H���   H�L$0���   H��(���������̉T$H�L$H��(H�4m H���   �T$8H�L$0���   H��(������������������H�L$H��(H��l H���   H�L$0���  H��(����������H�L$H��(H��l H���   H�L$0���   H��(���������̉T$H�L$H��(H��l H���   �T$8H�L$0��X  H��(������������������H��(H�]l H���   �PH��(�������H�L$H��(H�8l H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H��k H���   H�L$0���  H��(����������H�L$H��(H��k H���   H�L$0���  H��(����������L�L$ L�D$H�T$H�L$H��8H��k H���   H�L$hH�L$(�L$`�L$ L�L$XL�D$PH�T$HH�L$@���  H��8����������D�L$ L�D$H�T$H�L$H��(H�)k H���   D�L$HL�D$@H�T$8H�L$0���  H��(������������D�L$ L�D$H�T$H�L$H��8H��j H���   H�L$`H�L$ D�L$XL�D$PH�T$HH�L$@��   H��8������������������L�L$ L�D$H�T$H�L$H��(H�yj H���   L�L$HL�D$@H�T$8H�L$0��@  H��(������������D�L$ D�D$H�T$H�L$H��8H�)j H���   �L$h�L$(�L$`�L$ D�L$XD�D$PH�T$HH�L$@���  H��8������������H�L$H��(H��i H���   H�L$0���  H��(����������H�T$H�L$H��(H��i H���   H�T$8H�L$0���  H��(���������������̉T$H�L$H��(H�di H���   �T$8H�L$0���  H��(������������������L�D$H�T$H�L$H��(H�i H���   L�D$@H�T$8H�L$0���  H��(����������������������D�D$H�T$H�L$H��(H��h H���   D�D$@H�T$8H�L$0���  H��(����������������������D�D$H�T$H�L$H��(H�~h H���   D�D$@H�T$8H�L$0��   H��(����������������������D�D$H�T$H�L$H��(H�.h H���   D�D$@H�T$8H�L$0��  H��(����������������������H�T$H�L$H��(H��g H���   H�T$8H�L$0��  H��(����������������H�L$H��(H��g H���   H�L$0��  H��(�����������\$ D�D$H�T$H�L$H��hH�D$pH�L$xH�HH�D$pH��$�   H�HH�Ig H���   H��  H�L$XH��  H�L$PH�k  H�L$HH�/  H�L$@H�L$pH�IH�L$8H��$�   H�L$0��$�   �L$(��$�   �L$ ��$�   D��$�   H�L$pH�QH�L$p��  H��h����������������H��(H��f H�@��0  H��(�������H��(H�}f H�@��8  H��(�������H�L$H��(H�Xf H�@H�L$0��H  H��(�������������H�L$H��(H�(f H�@H�L$0��   H��(�������������H�L$H��(H��e H�@H�L$0��(  H��(�������������H�L$H��(H��e H�@H�L$0H�	��@  H�D$0H�     H��(��������������L�D$�T$H�L$H��H����H�D$0H�|$0 u3��^H�ie H�@H�D$     L�L$`D�D$XH�T$PH�L$0���  ��u'H�|$0 tH�/e H���   H�L$0�P H�D$0    H�D$0H��H����������������������L�L$ D�D$H�T$H�L$H��H�    �L$`�  H��d H�IH�L$0H�D$     L�L$hD��H�T$XH�L$PH�D$0���  H��H����������������D�L$ D�D$H�T$H�L$H��(H�id H�@D�L$HD�D$@H�T$8H�L$0��P  H��(���������������H�T$H�L$H��(H�#d H���   H�T$8H�L$0���  H��(����������������L�L$ L�D$H�T$H�L$H��HH��c H�@H��$�   H�L$0�L$x�L$(H�L$XH�L$ L�L$pL�D$hH�T$`H�L$P��X  H��H����������������H�L$H��xH�D$0����H�L$8�d  �H�L$(�i  �H��$�    tH�L$(��  H��u#�D$    H�L$(�  �H�L$8�Q����D$ �hH�L$(�  A�   H��H��$�   �����H�L$(�  H�D$XH��$�   H�D$8H�T$8�=��耣���D$$H�L$(�2  �H�L$8�����D$$H��x���������������H�L$H��xH�D$0����H�L$8�  �H�L$(�  �H��$�    tH�L$(�  H��u#�D$    H�L$(�  �H�L$8�q����D$ �hH�L$(��  A�   H��H��$�   �����H�L$(�  H�D$XH��$�   H�D$8H�T$8�<��蠢���D$$H�L$(�R  �H�L$8�����D$$H��x���������������D�D$�T$H�L$H��(H��a H���   D�D$@�T$8H�L$0���  H��(��������H�T$H�L$H��(H�sa H���   H�T$8H�L$0���  H��(����������������H��(H�=a H���   ��(  H��(��������������������H��(H�a H���   ���  H��(��������������������H�L$H��(H�D$0H� H�L$0�H��(��������������������H�T$H�L$H��(H�D$0H� H�T$8H�L$0�PH��(���������L�D$H�T$H�L$H��(H�D$0H� L�D$@H�T$8H�L$0�PH��(���������������L�L$ L�D$H�T$H�L$H��8H�D$@H� �L$`�L$ L�L$XL�D$PH�T$HH�L$@�PH��8�������������H�L$H��(��  H�L$0H�H�D$0H��(�H�T$H�L$H��(H�D$0�     H�D$0H�@    H��_ H��  H�T$8H�L$0�PXH�D$0H��(������H�T$H�L$H��(H�D$0�     H�D$0H�@    H�[_ H��  H�T$8H�L$0�PPH�D$0H��(�������L$H�L$H�D$�    H�D$�D$�@H�D$�����H�L$H�D$H�     H�D$H�@    H�D$H�@    H�D$�@    H�D$�@    H�D$H�@(    H�D$H�@     H�D$��������������H�L$H��(H�D$0H�������H�D$0H�     H��(����������H�L$H�D$H� ��̉T$�L$�D$�L$ȋ������������̉T$�L$�D$�L$ȋ�������������H��(H�^ H��  ��  H��(����L�L$ D�D$H�T$H�L$H��(H��] H��  L�L$HD�D$@H�T$8H�L$0�PH��(���������������H�L$H��(H��] H��  H�L$0���   H��(���������̉T$H�L$H��(H�d] H��  �T$8H�L$0��(  H��(��H�L$H��(H�8] H��  H�L$0���   H��(����������H�L$H��(H�] H��  H�L$0�PxH��(�������������H�L$H��(H��\ H��  H�L$0���   H��(����������H�T$H�L$H��(H��\ H��  H�T$8H�L$0�PxH��(���H�L$H��(H�x\ H���   H�L$0�PHH��(������������̉L$H��(H�I\ H���   3ҋL$0�H��(��������������H�L$H��(H�\ H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H��[ H���   H�L$0�PH��(�������������H�L$H��(H��[ H���   H�L$0�PH��(�������������H�L$H��(H�x[ H���   H�L$0�PPH��(�������������H�L$H��(H�H[ H���   H�L$0�PH��(������������̉T$�L$H��(H�[ H���   �T$8�L$0�H��(��������H�L$H��(H��Z H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H��Z H���   H�L$0�PPH��(�������������H�L$H��(H�xZ H���   H�L$0�PH��(�������������H�L$H��(H�HZ H���   H�L$0�PPH��(�������������H�L$H��(H�Z H���   H�L$0�PH��(������������̉L$H��(H��Y H���   �T$0�2  �H��(�����������H�L$H��(H��Y H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H�xY H���   H�L$0�PPH��(�������������H�L$H��(H�HY H���   H�L$0�PH��(�������������H�L$H��(H�Y H���   H�L$0�PPH��(�������������H�L$H��(H��X H���   H�L$0�PH��(�������������H�L$H��(H��X H���   H�L$0�PPH��(�������������H�L$H��(H��X H���   H�L$0�PH��(�������������H�L$H��(H�XX H���   H�L$0�P H��(������������̉L$H��(H�)X H���   3ҋL$0�H��(��������������H�L$H��(H��W H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H��W H���   H�L$0�PPH��(�������������H�L$H��(H��W H���   H�L$0�PH��(������������̉L$H��(H�YW H���   �T$0�'  �H��(�����������H�L$H��(H�(W H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H��V H���   H�L$0�PPH��(�������������H�L$H��(H��V H���   H�L$0�PH��(������������̉L$H��(H��V H���   �T$0�O  �H��(�����������H�L$H��(H�XV H���   H�L$0H�	�P H�D$0H�     H��(��������������H�T$H�L$VWH��HH�V H���   H�T$`H�L$ �H�|$hH��   �H�D$hH��H_^������������H�T$H�L$VWH��HH��U H���   H�T$`H�L$ �PH�|$hH��   �H�D$hH��H_^�����������H�T$H�L$VWH��HH�qU H���   H�T$`H�L$ �PH�|$hH��   �H�D$hH��H_^�����������H�T$H�L$VWH��   H�U H���   H��$�   H�L$ �PH��$�   H��`   �H��$�   H�Ĉ   _^������������H�T$H�L$H��(H��T H���   H�T$8H�L$0�P H��(�������������������H�T$H�L$H��(H��T H���   H�T$8H�L$0�P(H��(�������������������H�T$H�L$H��(H�CT H���   H�T$8H�L$0�P0H��(�������������������H�T$H�L$H��(H�T H���   H�T$8H�L$0�P8H��(������������������̉T$H�L$H��(H��S H���   �T$8H�L$0�PHH��(���������������������H�T$H�L$H��(H��S H���   H�T$8H�L$0�P@H��(�������������������H��(H�MS H���   3ҹ�  �H��(�����������������H�L$H��(H�S H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��(H��R H���   H�L$0�PPH��(�������������H�L$H��(H��R H���   H�L$0�PH��(�������������D�D$H�T$H�L$H��(H�nR H���   D�D$@H�T$8H�L$0�P(H��(��������̉L$H��(H�9R H���   3ҹ:  �H��(�������������H�L$H��(H�R H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H��8H�L$ �  �D$     H�D$(    L�D$ �   H�L$@�X0����u3��H�D$(H��8�������H��(H�}Q H���   3ҹ�F �H��(�����������������H�L$H��(H�HQ H���   H�L$0H�	�P H�D$0H�     H��(��������������H�T$H�L$H��8H�|$H u3��=H�L$ �   �D$     H�D$HH�D$(L�D$ �   H�L$@�/����u3���   H��8���������������������H��(H��P H���   3ҹ�_ �H��(�����������������H�L$H��(H�hP H���   H�L$0H�	�P H�D$0H�     H��(��������������H�L$H�D$�     H�D$H�@    H�D$��������������H�L$H��(H��O H���   H�L$0�PH��(�������������H�L$H��(H��O H���   H�L$0�PH��(������������̉T$H�L$H��(H��O H���   �T$8H�L$0�P H��(���������������������D�D$�T$H�L$H��(H�OO H���   D�D$@�T$8H�L$0�P(H��(����������̉T$H�L$H��(H�O H���   �T$8H�L$0�P0H��(���������������������H�L$H��(H��N H���   H�L$0�P8H��(������������̉T$H�L$H��(H��N H���   �T$8H�L$0�P@H��(���������������������D�D$�T$H�L$H��(H�_N H���   D�D$@�T$8H�L$0�PHH��(�����������L�L$ D�D$�T$H�L$H��8H�N H���   H�L$`H�L$ L�L$XD�D$P�T$HH�L$@���   H��8��������������������H�T$H�L$H��(H��M H���   H�T$8H�L$0�P`H��(�������������������H�T$H�L$H��(H��M H���   H�T$8H�L$0���   H��(����������������H�T$H�L$H��(H�CM H���   H�T$8H�L$0���   H��(����������������H�T$H�L$H��(H�M H���   H�T$8H�L$0���   H��(����������������H�L$H��(H��L H���   H�L$0�PhH��(�������������D�D$H�T$H�L$H��(H��L H���   D�D$@H�T$8H�L$0�PpH��(��������̉T$H�L$H��(H�TL H���   �T$8H�L$0�PxH��(���������������������H�T$H�L$H��H3�H�L$X�V���H�L$P�,����D$4�T$4H�L$X�:����D$0    �
�D$0���D$0�D$49D$0}AH�D$<H�D$ L�L$8A�����T$0H�L$P�y����T$8H�L$X������T$<H�L$X������H��H�������H�T$H�L$H��HH�T$,H�L$X�s����|$, ��   H�L$P�n���H�T$(H�L$X�O����|$( td�D$$    �
�D$$���D$$�D$(9D$$}FH�T$ H�L$X����H�T$0H�L$X�����
�D$ ���D$ �D$09D$ �T$ H�L$P�8�����릸   H��H�����������H��(H��J H���   �H��(��������H�L$H��(H��J H���   H�L$0H�	�PH�D$0H�     H��(��������������L�L$ L�D$H�T$�L$H��H  H��H H3�H��$0  �    �YJ �t  ��t�  �EJ �   �   �����   ������D$ ��$P  �J �4  �L$ �ы��'  ��u��   H��$p  H�D$(L�L$(L��$X  ��  H�L$0��� �   ��$P  ��  ��tH�x� �#  �!�   ��$P  ��  ��tH�e� �   H�L$0��  �   @��$P  �  ��tH��$h  H��$`  �   �    ��$P  �k  ��uH�� �  H�D$(    H��$0  H3��"R  H��H  �����������H��8�V� ��t
�D$    ��D$     �D$ H��8�������H�L$H��(H�L$0��� H��(��������H�L$H��(H�L$0��� H��(��������H�T$H�L$H��  H��F H3�H��$�  H�L$8����H�L$8����H�D$0L�L$0L��� �?   H�L$@�8� H��$�  H�D$(H��$�  H�D$ L�L$@L�Ҳ ��  H��$�   �   H��$�   �s   H��$�  H3���P  H�Ę  �����������̉T$�L$�D$�L$#ȋ�������������H��(�   �   �=���   ���1���    ���%��H��(�H�L$H��(H�T$0H��� �Ɠ��H��(��L�D$H�T$H�L$L�L$ H��HH�|$X 3���   H�D$hH�D$(L�L$(L�D$`H�T$XH�L$P�� H�H�D$ H�|$  |H�D$XH9D$ ��   H�|$  }^H�� �N  L�s� H�t� H������H�D$0�   @�   �X��L�ѱ A�2   H�L$0H�ы�������F ��t�H�D$XH�L$PH�H���@� H�D$XH��H�D$ H�D$(    H�D$ H��H�������������H�L$H�D$H�     H�D$H�@    H�D$�@    H�D$�@    H�D$���������������������H�L$H��(H�L$0�=  H��(���������H�T$H�L$H��(H�D$0H�     H�D$0H�@    H�D$0�@    H�D$0�@    H�D$8H�L$8�I9H��   A�   �   H�L$0��  ��u�  �   Hk� H�L$0H�	H�T$8���   Hk�H�L$0H�	H�T$8�R��   Hk�H�L$0H�	H�T$8�R��   Hk� H�L$0H�I�   �   A�   �   H�L$0�7  ��u�   �   Hk� H�L$0H�	H�T$8���   Hk�H�L$0H�	H�T$8�R��   Hk�H�L$0H�	H�T$8�R��   Hk�H�L$0H�	H�T$8�R��   Hk� H�L$0H�I�   H�D$0H��(�������������H�T$H�L$H��(H�D$0H�     H�D$0H�@    H�D$0�@    H�D$0�@    H�T$8H�L$0�  H�D$0H��(���������H�T$H�L$H��(H�T$8H�L$0�c  H�D$0H��(����������D�D$�T$H�L$H��8H�L$@��   �|$H ��   HcD$HH��H�aC H�IH�L$ L��� �I   ��H�D$ ���  H�L$@H�H�D$@H�8 u3��   �|$P tXHcD$PH��H�C H�IH�L$(L��� �N   ��H�D$(���  H�L$@H�AH�D$@H�x uH�D$@H��袐��3��!H�D$@�L$H�HH�D$@�L$P�H�   �3�H��8���������H�L$H��(H�D$0H���Z���H�D$0H��H���I���H�D$0�@    H�D$0�@    H��(�������������H�T$H�L$H��8H�L$@����H�|$H �H  H�D$HH�8 �9  H�D$H�x �*  H�D$HHc@H��H��A H�IH�L$ L��� �l   ��H�D$ ��P  H�L$@H�H�D$@H�8 u3���   H�D$HH�x tdH�D$H�x tYH�D$HHc@H��H��A H�IH�L$(L�{� �q   ��H�D$(��P  H�L$@H�AH�D$@H�x uH�L$@����3��oH�D$@H�L$H�I�HH�D$@H�L$H�I�HH�D$@D�@H�D$@H�H�D$HH��"  H�D$@H�x t H�D$@D�@H�D$@H�PH�D$HH�H�t"  �   H��8�����������L�L$ D�D$�T$H�L$H��HH�L$P����H�|$h ��  �|$X ��  HcD$XH��H��@ H�IH�L$ L��� ��   ��H�D$ ��P  H�L$PH�H�D$PH�8 u3��E  H�|$p tm�|$` tfHcD$`H��H�%@ H�IH�L$(L�u� ��   ��H�D$(��P  H�L$PH�AH�D$PH�x uH�L$P�L���3���   H�D$P�L$`�H�eH�D$P�@   H�D$PHc@H��H��? H�IH�L$0L�/� ��   ��H�D$0��P  H�L$PH�AH�D$PH�x uH�L$P�����3��kH�D$P�L$X�HH�D$PD�@H�D$PH�H�L$h��   H�|$p tH�D$PD�@H�D$PH�PH�L$p�   ��   Hk� H�L$PH�I�T$X��   H��H�������������������H�L$H�D$H�     H�D$H�@    H�D$�@    H�D$�@    ����������L�L$ L�D$�T$H�L$VWH���  W��D$(�D$$    3�H�L$`�4��3�H�L$H�4��3�H��$�   ��3��Hc�$�  H��$�  H�I�<�}W��[  ��$�   �C  H�L$0�jk��3�H��$�   �3���   Hk� H��$�  H�	HcHk�H�L$`H��$   H��H�4�   �   Hk�H��$�  H�	HcHk�H��$   H�H��L�D$`H��H��$�  �A��H��$�   H��H��   ��D$    �
�D$ ���D$ �   Hk� H��$�  H�I�9D$ ��   HcD$ H��$�  H�	Hc�Hk�H��$   H�H��L�D$`H��H��$�   �'A��H�L$HH��H��   �L�D$HH��$�   H��$0  �B��H��H�L$0��   H��$�   H�L$HH��H��   ��A���W�H��$�   蟾��H��$�   H��$  H��   �H�T$0H��$   �9��H��$  H�yHH��   ��D$0�2�����$�   �D$8������$�   f/���   �D$0� �����$�   �D$@������$�   f/���   H��$  H��HH��$�   W��҅ W�H��$`  �i��H��$�   L��H��H��$�  ��@��H��$  H�yH��   �H��$  H��H��$  H��HL��H��H��$�  �@��H��$  H�y0H��   ��S  �D$8�(����D$x�D$@�����L$xf/���   �� W�W�H��$P  �Ph��H��$  H��HL��H��H��$   �-@��H��$  H�yH��   �H��$  H��H��$  H��HL��H��H��$  ��?��H��$  H�y0H��   ��   W�W��{� H��$H  �g��H��$  H��HL��H��H��$x  �?��H��$  H�y0H��   �H��$  H��HH��$  H��0L��H��H��$�  �V?��H��$  H�yH��   �H��$  H��$h  �/��H��$  H��`   ��D$     �
�D$ ���D$ ��$�  9D$ }"HcD$ H��$�  H�I���L$$ȋ��D$$��HcD$$H��$�  H�	Hc�Hk�H��$   H�H��L��H��$  H��$�  �H  H�L$`H��H��   �D$$��H�H��$�  H�	Hc�Hk�H��$   H�H��L��H��$  H��$  ��  H�L$HH��H��   ��D$     �
�D$ ���D$ Hc�$�  H��$�  H�I��9D$ ��   �D$ ��Hc�$�  H��$�  H�RH��$�   �H��$�   �<��L$$ȋ�H�H��$�  H�	Hc�Hk�H��$   H�H��L��H��$  H��$8  �:  H��$�   H��H��   �L��$�   H�T$HH�L$`��  �L$(�X�(��D$(H�D$`H�L$HH��H��   �H�D$HH��$�   H��H��   �������D$(H���  _^����������������������L�L$ L�D$H�T$H�L$H��8H�D$@H�����H�Hk�H�L$HH�H��H�D$(H�L$@�[  �D$ �|$ �t!�|$  t2�|$ tJ�|$ tc�|$ t|�   H�D$P� ���H�D$X� ����|H�D$PH�L$(�	�H�D$XH�L$(�I��]H�D$PH�L$(�I�H�D$XH�L$(�I��=H�D$PH�L$(�I�H�D$XH�L$(�I��H�D$PH�L$(�I�H�D$XH�L$(�	�H��8�������D�D$�T$H�L$H��8H�L$@����D$$H�L$@�f  �D$ �D$$9D$Ht
�|$H���u�D$ 9D$Pt
�|$P���u�o�|$P���t�D$P�D$ �|$H���t�D$H�D$$�|$ �t#�D$ �L$$��H�L$@�	��   ��H�L$@��!�D$$����H�L$@�	��   ��H�L$@�H��8���������������������L�L$ L�D$H�T$H�L$H���   H�L$@��b���D$     �
�D$ ���D$ H��$   �@9D$ ��  HcD$ H��$   H�	H��H���&����u�HcD$ H��$   H�	H��H������H�Hk�H��$  H�H��H�D$(H�D$(H�L$(�I9H��   H�D$(Hc Hk�H��$  H�H��H�L$(HcIHk�H��$  H�H��L��H��H�L$X��8��H�D$0H�L$(Hc	Hk�H��$  H�H��H�T$(HcRHk�L��$  L�I��L��H��$�   �8��H�L$0L��H��H��$�   �9��H��H�L$@�  �   H�D$(Hc Hk�H��$  H�H��H�L$(HcIHk�H��$  H�H��L��H��H�L$p�'8��H�D$8H�L$(HcIHk�H��$  H�H��H�T$(HcRHk�L��$  L�I��L��H��$�   ��7��H�L$8L��H��H��$�   ��8��H��H�L$@��  ����H�T$@H��$  � 0��H��$  H���   �����������������L�L$ L�D$H�T$H�L$H��xH�L$0�  �D$     �
�D$ ���D$ H��$�   �@9D$ �  HcD$ H��$�   H�	H��H��������u�HcD$ H��$�   H�	H��H���g��H�Hk�H��$�   H�H��H�D$(H�D$(Hc Hk�H��$�   H�H��H��H�L$0�7  H�D$(Hc@Hk�H��$�   H�H��H��H�L$0�  H�D$(Hc@Hk�H��$�   H�H��H��H�L$0��  H�D$(H�L$(�I9Ht(H�D$(Hc@Hk�H��$�   H�H��H��H�L$0�  �����L��$�   H��$�   H�L$0�  H��x����������H�L$H��8�D$$    H�D$@�x|H�D$@H�8 u3��O�D$     �
�D$ ���D$ H�D$@�@9D$ })HcD$ H�L$@H�	H��H���  ��t
�D$$���D$$뿋D$$H��8�����������������̉T$H�L$H��8�D$H�D$ �
�D$ ���D$ H�D$@�@9D$ }/HcD$ H�L$@H�	H��H���(  ��t�D$H�L$ +ȋ����빸����H��8��������̉T$H�L$H��8�|$H |H�D$@H�8 u������N�D$     �
�D$ ���D$ H�D$@�@9D$ }'HcD$ H�L$@H�	H��H���
��;D$Hu�D$ ��������H��8�������̉T$H�L$H��8�D$  �D$$    �
�D$$���D$$H�D$@�@9D$$}OHcD$$H�L$@H�	H��H���	��;D$Hu.�D$ �D$(HcL$$H�T$@H�H���.  ���L$(ȋ��D$ ��D$ ��H��8������������������H�L$H��8�D$$    �D$     �
�D$ ���D$ H�D$@�@9D$ }*HcD$ H�L$@H�	H��H���d  ���t
�D$$���D$$뾋D$$H��8�����������H�L$H��8�D$$    �D$     �
�D$ ���D$ H�D$@�@9D$ })HcD$ H�L$@H�	H��H��������t
�D$$���D$$뿋D$$H��8������������H�L$H��8�D$     �
�D$ ���D$ H�D$@�@9D$ }&HcD$ H�L$@H�	����HcL$ H�T$@H������D$     �
�D$ ���D$ H�D$@�@9D$ ��   HcD$ H�L$@H�	��%   �����   HcD$ H�L$@H�	H��H�������D$(�D$ ���D$$�
�D$$���D$$H�D$@�@9D$$}EHcD$$H�L$@H�	H��H�����;D$(u$HcD$$H�L$@H�	����HcL$$H�T$@H�����<���H��8�������������H��8�   �  H�D$ H�|$  u3��H�D$ �PH��8���������������������H�L$H��8H�D$@H�8 u�?�   ��  H�D$ H�|$  u�&H�D$@H� H�D$(H�L$(H�D$ �PH�D$@H�     H��8�������H�T$H�L$H��8�   �h  H�D$ H�|$  tH�D$ H�x u3��H�T$HH�L$@H�D$ �PH��8���������������������H�T$H�L$H��8�    �  H�D$ H�|$  tH�D$ H�x  u3��H�T$HH�L$@H�D$ �P H��8���������������������D�L$ D�D$H�T$H�L$H��8�(   �  H�D$ H�|$  tH�D$ H�x( u3��D�L$XD�D$PH�T$HH�L$@H�D$ �P(H��8�����������������H�T$H�L$H��8�0   �8  H�D$ H�|$  tH�D$ H�x0 u3��H�T$HH�L$@H�D$ �P0H��8���������������������H�T$H�L$H��8�8   ��  H�D$ H�|$  tH�D$ H�x8 u3��H�T$HH�L$@H�D$ �P8H��8��������������������̉T$H�L$H��8�@   �y  H�D$ H�|$  tH�D$ H�x@ u2���T$HH�L$@H�D$ �P@H��8�������H�L$H��8�H   �-  H�D$ H�|$  tH�D$ H�xH u3��H�L$@H�D$ �PHH��8���������������H�L$H��8�P   ��  H�D$ H�|$  tH�D$ H�xP u3��H�L$@H�D$ �PPH��8��������������̉T$H�L$H��8�X   �  H�D$ H�|$  tH�D$ H�xX u3���T$HH�L$@H�D$ �PXH��8�������D�D$�T$H�L$H��8�`   �4  H�D$ H�|$  tH�D$ H�x` u������D�D$P�T$HH�L$@H�D$ �P`H��8����������H�L$H��8�h   ��
  H�D$ H�|$  tH�D$ H�xh u3��H�L$@H�D$ �PhH��8���������������H�T$H�L$H��8�p   �
  H�D$ H�|$  tH�D$ H�xp u�H�T$HH�L$@H�D$ �PpH��8�������H�T$H�L$H��8�x   �8
  H�D$ H�|$  tH�D$ H�xx u�H�T$HH�L$@H�D$ �PxH��8�������H�T$H�L$H��8��   ��	  H�D$ H�|$  tH�D$ H���    u3��H�T$HH�L$@H�D$ ���   H��8��������������̉T$H�L$H��8��   �	  H�D$ H�|$  tH�D$ H���    u��T$HH�L$@H�D$ ���   H��8�������������������H�L$H��8��   �-	  H�D$ H�|$  tH�D$ H���    u3��H�L$@H�D$ ���   H��8���������H�L$H��8��   ��  H�D$ H�|$  tH�D$ H���    u3��H�L$@H�D$ ���   H��8���������H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u�H�L$@H�D$ ���   H��8�����������H�L$H��8��   �=  H�D$ H�|$  tH�D$ H���    u�H�L$@H�D$ ���   H��8�����������H�L$H��8��   ��  H�D$ H�|$  tH�D$ H���    u�H�L$@H�D$ ���   H��8�����������D�D$�T$H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u3��D�D$P�T$HH�L$@H�D$ ���   H��8�������D�D$H�T$H�L$H��8��   �3  H�D$ H�|$  tH�D$ H���    u3��D�D$PH�T$HH�L$@H�D$ ���   H��8���������������������L�L$ L�D$�T$H�L$H��H��   �  H�D$0H�|$0 tH�D$0H���    u�2H�D$xH�D$(H�D$pH�D$ L�L$hL�D$`�T$XH�L$PH�D$0���   H��H�����������D�L$ L�D$�T$H�L$H��8��   �?  H�D$ H�|$  tH�D$ H���    u3��D�L$XL�D$P�T$HH�L$@H�D$ ���   H��8�������������D�D$H�T$H�L$H��8��   ��  H�D$ H�|$  tH�D$ H���    u3��D�D$PH�T$HH�L$@H�D$ ���   H��8���������������������D�D$�T$H�L$H��8��   �d  H�D$ H�|$  tH�D$ H���    u3��D�D$P�T$HH�L$@H�D$ ���   H��8�������L�D$H�T$H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u3��L�D$PH�T$HH�L$@H�D$ ���   H��8���������������������H�T$H�L$H��8��   �  H�D$ H�|$  tH�D$ H���    u3��H�T$HH�L$@H�D$ ���   H��8���������������L�D$H�T$H�L$H��8��   �3  H�D$ H�|$  tH�D$ H���    u3��L�D$PH�T$HH�L$@H�D$ ���   H��8���������������������D�L$ L�D$H�T$H�L$H��X�   �  H�D$@H�|$@ tH�D$@H��    u������DH��$�   H�D$0H��$�   H�D$(��$�   �D$ D�L$xL�D$pH�T$hH�L$`H�D$@��   H��X�������������������D�L$ L�D$H�T$H�L$H��X�  �  H�D$@H�|$@ tH�D$@H��   u������DH��$�   H�D$0H��$�   H�D$(��$�   �D$ D�L$xL�D$pH�T$hH�L$`H�D$@��  H��X�������������������D�L$ D�D$H�T$H�L$H��H�  �~  H�D$0H�|$0 tH�D$0H��   u3��)H�D$pH�D$ D�L$hD�D$`H�T$XH�L$PH�D$0��  H��H����������������̉T$H�L$H��8�  �	  H�D$ H�|$  tH�D$ H��   u3���T$HH�L$@H�D$ ��  H��8�����������������H�T$H�L$H��8�   �  H�D$ H�|$  tH�D$ H��    u�H�T$HH�L$@H�D$ ��   H��8�����������������L�D$�T$H�L$H��8�(  �D  H�D$ H�|$  tH�D$ H��(   u3��L�D$P�T$HH�L$@H�D$ ��(  H��8�������D�L$ L�D$�T$H�L$H��8�0  ��   H�D$ H�|$  tH�D$ H��0   u3��D�L$XL�D$P�T$HH�L$@H�D$ ��0  H��8�������������L�D$H�T$H�L$H�D$H�L$�@�\AH�D$��Y�(�H�D$H�L$�H�\IH�D$��Y�(��X�H�D$H�L$�H�\IH�D$��Y�(��X�������������̉L$H��(L�� �T$0�_� �  H��(���������������D�D$H�T$H�L$H��(HcD$@H��L��H�T$0H�L$8�&  H��(��������������H�L$VWH��XH�D$pH���`K��H�D$pH��H���OK����z H�L$ ����H�D$ H�|$pH��   ���z H�L$8迟��H�D$pH�L$8H�xH��   �H�D$p�@0    H�D$pH��X_^�����������������T$H�T$H�L$H��8H�D$H�@�YD$PH�D$H�H�YL$PH�D$H��YT$P�T$ (�(��D$ (�H�L$@�bJ��H�D$@H��8�����L�D$H�T$H�L$H��8H�D$HH�L$P�@(�YH�D$H�H�X�(�H�D$HH�L$P�H@�YI�X�H�D$HH�L$P�HX�YI�X�H�D$HH�L$P�H �Y	H�D$H�P�X�(�H�D$HH�L$P�P8�YQ�X�H�D$HH�L$P�PP�YQ�X�H�D$HH�L$P�P�YH�D$H��X�(�H�D$HH�L$P�X0�YY�X�H�D$HH�L$P�XH�YY�X��T$ (�(��D$ (�H�L$@�'I��H�D$@H��8����������H�T$H�L$H�D$H�L$� �XH�D$� H�D$H�L$�@�XAH�D$�@H�D$H�L$�@�XAH�D$�@H�D$����������H�T$H�L$VWH�D$�x0 ��   H�D$H�L$ � f/vH�D$H�L$ �� H�D$H�L$ �@f/AvH�D$H�L$ �A�@H�D$H�L$ �@f/AvH�D$H�L$ �A�@H�D$ H�L$� f/AvH�D$H�L$ ��@H�D$ H�L$�@f/A vH�D$H�L$ �A�@ H�D$ H�L$�@f/A(vH�D$H�L$ �A�@(�6H�D$H�xH�t$ �   �H�D$H�|$H�p�   �H�D$�@0   _^�����H�L$H�D$� %   @��t������H�D$� %���3ҹ   ����������������L�D$H�T$H�L$VWH��   H��$�   �x0 ��   H��$�   H��H��$�   L��H��H�L$8�"����~ H��H�L$P�����H��$�   H��   �H��$�   H��L��$�   H��H�L$h�Z��H��$�   H��   ��;W�H�L$ ����H�D$ H��$�   H��   �H��$�   H��$�   �   �H�Ĉ   _^��H�L$H�D$� %    ���������������H�L$H��8H�L$@�����D$ �|$ �u3���D$ �   �L$$�ȋD$$��H��8����H�T$H�L$H��(H�s H���   H�T$8H�L$0���   H��(����������������H�L$H��(H�D$0H�8 u�H�+ H���   H�L$0���   H��(�������������L�L$ L�D$H�T$H�L$H��8H�� H���   H�L$`H�L$ L�L$XL�D$PH�T$HH�L$@�H��8����������������������L�L$ L�D$H�T$H�L$H��8H�� H���   H�L$`H�L$ L�L$XL�D$PH�T$HH�L$@���  H��8������������������L�L$ L�D$H�T$H�L$H��(H�) H���   L�L$HL�D$@H�T$8H�L$0�PH��(���������������L�L$ L�D$H�T$H�L$H��8H�� H���   H�L$hH�L$(H�L$`H�L$ L�L$XL�D$PH�T$HH�L$@�P@H��8�����������D�D$�L$H�L$H��(H�} H���   D�D$@�L$8H�L$0��x  H��(��������������������D�D$�L$H�L$H��(H�- H���   D�D$@�L$8H�L$0���  H��(��������������������D�D$H�T$H�L$H��(H�� H���   D�D$@H�T$8H�L$0���  H��(����������������������D�D$H�T$H�L$H��(H�� H���   D�D$@H�T$8H�L$0���  H��(����������������������L�L$ L�D$H�T$H�L$VWH��hH�7 H���   H��$�   H�L$8H��$�   H�L$0��$�   �D$(��$�   �D$ L��$�   L��$�   H��$�   H�L$@���  H��$�   H��   �H��$�   H��h_^�������������L�L$ L�D$H�T$H�L$VWH��hH�� H���   H��$�   H�L$0��$�   �D$(��$�   �D$ L��$�   L��$�   H��$�   H�L$@���  H��$�   H��   �H��$�   H��h_^����������D�D$H�T$H�L$H��hH�D$(�����D$     H�L$@袕�����$�   H�L$0�@:��H��H�L$P�3#���E3�L�D$@H�T$PH�L$p�����H�L$P�$��H�T$@H�L$x�Q����D$ ���D$ H�L$@�<���H�D$xH��h�������������������L�L$ L�D$H�T$H�L$H��8H�9 H���   H�L$`H�L$ L�L$XL�D$PH�T$HH�L$@��   H��8�����������������̉T$H�L$H��(H�� H���   �T$8H�L$0��(  H��(������������������H��(H�� H���   ���   H��(��������������������H�L$H��(H�D$0H�8 u�H�k H���   H�L$0���   H��(�������������D�L$ D�D$H�T$H�L$H��XH�) H���   H��$�   H�L$@H��$�   H�L$8H��$�   H�L$0��$�   �L$(��$�   �L$ D�L$xD�D$pH�T$hH�L$`��P  H��X���������������D�L$ D�D$H�T$H�L$H��xH�� H���   H��$�   H�L$hH��$�   H�L$`H��$�   H�L$X��$�   �L$PH��$�   H�L$HH��$�   H�L$@H��$�   H�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ D��$�   D��$�   H��$�   H��$�   ���  H��x������������������D�L$ D�D$H�T$H�L$H��   H�� H���   H��$   H�L$pH��$�   H�L$hH��$�   H�L$`��$�   �L$XH��$�   H�L$PH��$�   H�L$HH��$�   H�L$@H��$�   H�L$8H��$�   H�L$0��$�   �L$(��$�   �L$ D��$�   D��$�   H��$�   H��$�   ���  H�Ĉ   �����������������L�L$ D�D$�T$H�L$H��HH�� H���   ��$�   �L$8��$�   �L$0�L$x�L$(H�L$pH�L$ L�L$hD�D$`�T$XH�L$P���   H��H����������������������L�L$ D�D$�T$H�L$H��HH�J H���   ��$�   �L$8��$�   �L$0�L$x�L$(H�L$pH�L$ L�L$hD�D$`�T$XH�L$P���   H��H����������������������D�D$�T$H�L$H��(H�� H���   D�D$@�T$8H�L$0���   H��(��������D�D$�T$H�L$H��(H�� H���   D�D$@�T$8H�L$0���   H��(��������D�D$�T$H�L$H��(H�O H���   D�D$@�T$8H�L$0���   H��(��������L�L$ L�D$H�T$H�L$H��HH�	 H���   ��$�   �L$8H��$�   H�L$0�L$x�L$(�L$p�L$ L�L$hL�D$`H�T$XH�L$P��0  H��H��������������������L�L$ L�D$H�T$H�L$H��HH�� H���   ��$�   �L$8H��$�   H�L$0�L$x�L$(�L$p�L$ L�L$hL�D$`H�T$XH�L$P��8  H��H��������������������L�L$ L�D$H�T$H�L$H��HH�	 H���   ��$�   �L$8H��$�   H�L$0�L$x�L$(�L$p�L$ L�L$hL�D$`H�T$XH�L$P��@  H��H��������������������D�L$ D�D$H�T$H�L$H��8H�� H���   �L$h�L$(H�L$`H�L$ D�L$XD�D$PH�T$HH�L$@��  H��8����������L�L$ D�D$H�T$H�L$H��8H�) H���   �L$`�L$ L�L$XD�D$PH�T$HH�L$@��  H��8��������������������D�L$ D�D$H�T$H�L$H��(H�� H���   D�L$HD�D$@H�T$8H�L$0���   H��(�����������̉T$H�L$H��(H�� H���   �T$8H�L$0���   H��(������������������D�L$ D�D$�T$H�L$H��8H�: H���   �L$`�L$ D�L$XD�D$P�T$HH�L$@��H  H��8����������������������D�L$ D�D$�T$H�L$H��(H��
 H���   D�L$HD�D$@�T$8H�L$0���   H��(��������������\$ �T$�L$H�L$H��8H��
 H���   H�L$`H�L$ �\$X�T$P�L$HH�L$@��   H��8������������D�L$ D�D$H�T$�L$H��(H�D$8�L$@�H�D$8�L$H�HL�D$8�   �L$0�S��H��(�����������D�D$�T$H�L$�   �������������L�D$�T$�L$H��8H�|$P tH�D$PH�8 t
H�D$PH� �f�   �L$@�S��H�D$(H�|$( u3��GH�L$(��R��H�D$ H�|$  u3��,H�|$P tH�D$PH�L$ H�H�D$ �@9D$H~3��H�D$ H��8�������̉T$H�L$H��HH�$	 H�@(�T$XH�L$P���   �D$ �|$  u3��   �D$ ��H�� H�IH�L$0L��u �	   ��H�D$0���  H�D$(H�|$( u3��G�D$ ��H�� H�I(H�L$8D�L$XD��H�T$(H�L$PH�D$8���   HcD$ H�L$(� H�D$(H��H�����������H�T$H�L$H��hH�� H3�H�D$P�D$,    �D$x�D$0�D$$    HcD$$�D@0�D$$���D$$HcD$$�D@x�D$$���D$$�D$(   ��D$(���D$(�|$( |X�D$(�ȋD$0�����D$ �D$ ��
}�D$ ��0HcL$$�D@�D$$���D$$��D$ ��7HcL$$�D@�D$$���D$$�HcD$$H�D$8H�|$8s��6  H�D$8�D@ E3�H�T$@H�L$p��4���D$,���D$,H�D$pH�L$PH3��m  H��h���������H�T$H�L$H��  HǄ$�   �����D$0    H��$�     @��   E3�H��s H��$�   �N4��H�D$xH�D$xH�D$PH��$�  H���H*��^�t f�D$(0 �D$     A�   E3�(�H��$   ��  H��$�   H��$�   H��$�   L�D$PH��$�   H��$�  �p����D$0���D$0H��$   ��3���H��$�   �3��H��$�  �S  ��  H��$�     ��   E3�H�s H��$�   �k3��H�D$`H�D$`H�D$pH��$�  H��
�H*��^�s f�D$(0 �D$     A�   E3�(�H��$P  ��  H��$�   H��$�   H��$�   L�D$pH��$�   H��$�  草���D$0���D$0H��$P  ��2���H��$�   ��2��H��$�  �p  ��   H��$�     ��   E3�H�-r H��$  �2��H��$�   H��$�   H��$�   �H*�$�  �^�r f�D$(0 �D$     A�   E3�(�H��$�   �
  H��$�   H��$�   H�D$8L��$�   H�T$8H��$�  諈���D$0���D$0H��$�   ��1���H��$  ��1��H��$�  �   E3�H�fq H��$h  �1��H�D$@H�D$@H�D$X��$�  H��$8  �1��H�D$HH�D$HH�D$hL�D$XH�T$hH��$�  �����D$0���D$0H��$8  �k1���H��$h  �]1��H��$�  H�Ĉ  �������������������H�L$H��(E3�A��  H�� H�L$0荨��H�� H��(������������������H�L$H��(E3�A��  H�� H�L$0�M���H�� H��(������������������H�L$H��(�� H�L$0�8  ��t$H�L$0�����E3�A��  H�J H�������H��o H�2 �{  H�& H��(������������������H�L$H��XH�D$0����H�T$8H�L$`�o��H�D$ H�D$ H�D$(E3�A��  H�� H�L$(�v����H�L$8��/��H�� H��X����������������H�L$H��XH�D$0����H�T$8H�L$`�o��H�D$ H�D$ H�D$(E3�A��  H�` H�L$(�����H�L$8�/��H�D H��X���������������̉T$H�L$H��(H�� H��  �T$8H�L$0�PH��(�����D�L$ D�D$�L$H�L$H��xH�D$H�����D$0    H�� H�@(��$�   f�L$(��$�   �L$ D��$�   D��$�   ��$�   H�L$P�PHH�D$8H�D$8H�D$@H�T$@H��$�   �a.���D$0���D$0H�L$P�.��H��$�   H��x���%8� ��������H�T$H�L$H�D$H��n H�H�D$��H�T$H�L$H�D$ÉT$H�L$H��(�D$8����tFL�o  H�D$0D�@��   H�L$0�9  �D$8����tH�D$0H��H����-��H�D$0H���$H�L$0�&  �D$8����t
H�L$0��-��H�D$0H��(����������H��8A��   L�'n �   �   �o� H�D$ H�L$ �� H��	 H��	 H��	 H�|$  u�   �+H�D$ H�     �  H��  �^  H�'  �R  3�H��8������������eH�%0   �������L�D$�T$H�L$H��   ��$�    u �=�  ~�� �ȉ� �3��`  ��$�   �(  H�D$H    ����H�@H�D$h�D$4    H�D$hH��$�   H�� 3�H��$�   �H�H�D$HH�|$H tH�D$hH9D$Hu
�D$4   �븋� ��t�   �  �E��    H�EB H�? �  ��t3��  H��= H�0; ��  �]    �|$4 u3�H�9 H�H�=f  t+H�] �  ��tL��$�   �   H��$�   �9 �   ��~ �d ���\ �%  ��$�    �  H�D$`    �_���H�@H�D$x�D$0    H�D$xH��$�   H�� 3�H��$�   �H�H�D$`H�|$` tH�D$xH9D$`u
�D$0   �븋| ��t�   �w  �  H�} ��| H�D$(H�|$( �[  H�G ��| H�D$ H�D$p    H�D$(H�D$8H�D$ H�D$@3�����   H�D$X    H�D$P    H�D$ H��H�D$ H�D$(H9D$ rH�D$ H�8 t3��}| H�L$ H9u��H�D$(H9D$ s�   H�D$ H��J| H�D$p3��E| H�L$ H��T$pH�� �$| H�D$XH�x �| H�D$PH�D$XH9D$8uH�D$PH9D$@t(H�D$XH�D$8H�D$8H�D$(H�D$PH�D$@H�D$@H�D$ �	���H�|$(�t�   H�L$(��| 3���{ H� H�� H� ��     �|$0 u3�H�� H��   H�Ę   ����������L�D$�T$H�L$H��(�|$8u�  L�D$@�T$8H�L$0�   H��(�����������L�D$�T$H�L$H��8�D$    �D$H��� �|$H u�=��  u�D$     �  �|$Ht�|$HuLH�=Ii  tL�D$P�T$HH�L$@�3i �D$ �|$  tL�D$P�T$HH�L$@�����D$ �|$  u�   L�D$P�T$HH�L$@�b(���D$ �|$HuE�|$  u>L�D$P3�H�L$@�?(��L�D$P3�H�L$@�.���H�=�h  tL�D$P3�H�L$@��h �|$H t�|$HuHL�D$P�T$HH�L$@�������u�D$     �|$  t"H�=fh  tL�D$P�T$HH�L$@�Ph �D$ ��D$     ��� �����D$ H��8���%X{ �%J{ �%<{ ������������H��HH�=�  t
H�=�  uOH�=�  u
H�=�  t;H�h H�D$(H��h H�D$ E3�A�E   H��h �   �Qz ��u�3�H�=�  t3��g�D$ M   L�i A�   �   �    �z H�D$0H�L$0��x H�W H�P H�1 H�|$0 u�   �H�D$0H�     3�H��H����������������H�L$H��HH� ��x H�D$ H�|$ �uH�L$P��y �   �   �o
  �H�� �Ux H�D$ H�� �Cx H�D$(H�L$P�;x L�D$(H�T$ H���E
  H�D$0H�L$ �x H�� H�L$(�x H�X �   � 
  H�D$0H��H�����H�L$H��8H�L$@�-���H��u
�D$ ������D$     �D$ H��8���%>y �%0y �%"y �%y ����L�L$ L�D$H�T$H�L$H��(H�D$HL�@8H�T$HH�L$8�   �   H��(�������L�D$H�T$H�L$H��XH�D$p� ����D$ H�D$`H�D$8H�D$p� ������t)H�D$pHc@H�L$`H�H��H�L$p�I��Hc�H#�H�D$8HcD$ H�L$8H�H�D$0H�D$hH�@�@H�L$hHAH�D$@H�D$`H�D$(H�D$@�@$����t&H�D$@�@��$��k�H�H�L$(H�H��H�D$(H�D$(H�L$0H3�H��H�D$0H�L$0�   H��X���������������ff�     H;)� uH��f����u��H���   ��%w �%�v �%�v �%�v �%�v �%�v �%�v �%�v �%�v �%�v ����H�L$H��(��u ��� �   ��  H�L$0��  �=��  u
�   ��  �	 ���  H��(������H�L$H��8�   ��  ��t�   �)H��� �  H�D$8H��� H�D$8H��H�B� H��� H�� H�D$@H�� ��� 	 ����    ���    �   Hk� H��� H�   �   Hk� H��� H�L �   Hk�H��� H�L H�e �����H��8����������������H��(�   �   H��(�������������̉L$H��(�   ��  ��t�D$0���)H��� �  H�D$(H��� H�D$(H��H�B� H��� H�� ��� 	 ����    ���    �   Hk� H��� �T$0H�H�7d ����H��(������L�D$�T$�L$H��8�   �A  ��t�D$@���)H�"� ��  H�D$8H�	� H�D$8H��H��� H��� H�c� �I� 	 ��C�    �|$H vH�|$P u�D$H    �|$Hv
�D$H�ȉD$H�D$H���#� �   Hk� H�� �T$@H��D$     �
�D$ ���D$ �D$H9D$ s"�D$ �L$ ����H��� L�D$PI��H����H�$c ����H��8��%�s ������������L�L$ D�D$H�T$H�L$H��8�D$     HcD$PH�L$HH��H��H�L$@H�H��H�D$@�D$P�ȉD$P�|$P | H�D$HH�L$@H+�H��H�D$@H�L$@�T$X���D$    �|$  uL�L$XD�D$PH�T$HH�L$@�F   H��8��H�L$H��8H�D$@H� H�D$(H�D$(� �D$ �|$ csm�t��F  3�H��8��������L�L$ D�D$H�T$H�L$H��8�D$P�ȉD$P�|$P | H�D$HH�L$@H+�H��H�D$@H�L$@�T$X��� H��8��%jr �%lr �%nr �%pr �%rr ��H�T$H�L$H��(H�D$0Hc@<H�L$0H�H��H�D$�$    H�D$�@H�L$H�DH�D$��$���$H�D$H��(H�D$H�D$�@9$s1H�D$�@H9D$8r H�D$�@H�L$A��H9D$8sH�D$��3�H��(�������������H�L$H��XH����H�D$0H�L$0�q   ��u3��bH�D$0H�L$`H+�H��H�D$@H�T$@H�L$0����H�D$8H�|$8 u3��-H�D$8�@$%   ���u
�D$    ��D$     �D$ �3�� H��X���H�L$H��(H�D$0H�$H�$� =MZ  t3��NH�$Hc@<H�$H�H��H�D$H�D$�8PE  t3��&H�D$H��H�D$H�D$� =  t3���   H��(����������H��HH�D$(    H�2��-�+  H9�� tH��� H��H��� ��   H�L$(��o H�D$(H�D$ �Oo ��H�L$ H3�H��H�D$ �?o ��H�L$ H3�H��H�D$ H�L$0�*o �D$0H�� H3D$0H�L$ H3�H��H�D$ H�D$ H�L$ H3�H��H�D$ H�������  H�L$ H#�H��H�D$ H�2��-�+  H9D$ uH�3��-�+  H�D$ H�D$ H��� H�D$ H��H��� H��H���������������H�\$WH�� H��q H�=�r H;�s H�H��t��H��H;�r�H�\$0H�� _���H�\$WH�� H��s H�=�t H;�s H�H��t��H��H;�r�H�\$0H�� _��%o �%�o ������H��(H�=� �T   H��(���%�n �%�n �% o �%o �%o �%o �%o �%o �%o �%o �%o �%o �%o �%o �%�m �%�m �%�m �%�m �%xm �%jm �%\m �%�m ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@UH�� H��H�Mh�YZ��H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H���   �&Z��H�� ]����������������������@UH�� H��L�8v  A�E   H��0 H�M ��Y��H�� ]���������������������@UH�� H��H�M@�Y��H�� ]�@UH�� H��E ����t�e �H�Mp�Y��H�� ]�������������������@UH�� H��H���   軗��H�� ]�@UH�� H��H���   蠗��H�� ]�@UH�� H��H���   �0Y��H�� ]�@UH�� H��H���   �Y��H�� ]�������������������������������������@UH�� H��H�MP��X��H�� ]�@UH�� H��H�Mh��X��H�� ]�����������������@UH�� H��H�M@����H�� ]�@UH�� H��L�Hu  A�;   H�#/ H�M(�YX��H�� ]�@UH�� H��H�M@�UX��H�� ]�@UH�� H��H�M`�=X��H�� ]�@UH�� H��E4����t�e4�H���   �X��H�� ]�@UH�� H��H�MH��W��H�� ]�@UH�� H��H�M`��W��H�� ]�@UH�� H��E4����t�e4�H���   �W��H�� ]�@UH�� H��H���   �W��H�� ]�@UH�� H��H�MH�W��H�� ]�@UH�� H��H�M`�pW��H�� ]�@UH�� H��E0����t�e0�H���   �GW��H�� ]�@UH�� H��H�Mx�/W��H�� ]�@UH�� H��H���   �W��H�� ]�@UH�� H��H�M@��V��H�� ]�@UH�� H��H�Mh��V��H�� ]�@UH�� H��E4����t�e4�H���   �V��H�� ]�@UH�� H��H���   �V��H�� ]�@UH�� H��H���   �V��H�� ]�@UH�� H��H���   �jV��H�� ]�@UH�� H��H���   �OV��H�� ]�@UH�� H��E ����t�e �H���   �&V��H�� ]�@UH�� H��E ����t�e �H���   ��U��H�� ]�@UH�� H��H���   ��U��H�� ]�@UH�� H��E ����t�e �H���   �U��H�� ]�@UH�� H��E ����t�e �H���   �U��H�� ]����������������@UH�� H��H�M@�iU��H�� ]�@UH�� H��E ����t�e �H�Mx�CU��H�� ]���@UH�� H��H�M@�~���H�� ]�@UH�� H��E ����t�e �H���   �U���H�� ]����������������@UH�� H��H�M@��T��H�� ]�@UH�� H��H�M@��T��H�� ]�@UH�� H��H�M@�T��H�� ]�@UH�� H��H�M@�T��H�� ]�@UH�� H��H�M@�yT��H�� ]�@UH�� H��H�M@�aT��H�� ]�@UH�� H��E ����t�e �H�Mx�;T��H�� ]�@UH�� H��H�M@�x���H�� ]�@UH�� H��E ����t�e �H���   �O���H�� ]�@UH�� H��H�M@�7���H�� ]�@UH�� H��E ����t�e �H���   ����H�� ]�@UH�� H��H�M@�����H�� ]�@UH�� H��E ����t�e �H���   �xS��H�� ]�@UH�� H��H�M0赑��H�� ]�@UH�� H��E ����t�e �H�Mp菑��H�� ]�@UH�� H��H�M@�"S��H�� ]�@UH�� H��E ����t�e �H�Mx��R��H�� ]�@UH�� H��H�M0��R��H�� ]�@UH�� H��H�MH��R��H�� ]�@UH�� H��H�M@�R��H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��E ����t�e �H���   �Ȑ��H�� ]�@UH�� H��H�M@谐��H�� ]�@UH�� H��E ����t�e �H���   臐��H�� ]�@UH�� H��H�M@�R��H�� ]�@UH�� H��E ����t�e �H�Mx��Q��H�� ]�@UH�� H��H�M8�1���H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��E ����t�e �H���   �����H�� ]�@UH�� H��H�M@�؏��H�� ]�@UH�� H��E ����t�e �H���   诏��H�� ]�@UH�� H��E ����t�e �H���   膏��H�� ]�@UH�� H��E ����t�e �H�M`�`���H�� ]�@UH�� H��E ����t�e �H���   �7���H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��E ����t�e �H���   �����H�� ]�@UH�� H��H�M@�P��H�� ]�@UH�� H��E ����t�e �H�Mp�cP��H�� ]���@UH�� H��H���   蛎��H�� ]�@UH�� H��H�Mp�.P��H�� ]�@UH�� H��H���   �h���H�� ]�@UH�� H��H��(  �M���H�� ]�@UH�� H��H��   �2���H�� ]�@UH�� H��H���   ����H�� ]��@UH�� H��H�M@�O��H�� ]�@UH�� H��E ����t�e �H�Mx�O��H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��H�M@���H�� ]�@UH�� H��E ����t�e �H�Mh���H�� ]�@UH�� H��H�M@H���F��H�� ]�@UH�� H��H�M@H���*��H�� ]�@UH�� H��L��r  A��   H�% H�M �N��H�� ]�@UH�� H��H�MH�O��H�� ]�@UH�� H��H�M`�N��H�� ]���������@UH�� H��H�Mh�nO��H�� ]�@UH�� H��H�M8�VO��H�� ]�@UH�� H��E0����t�e0�H���   � ��H�� ]�@UH�� H��H�M`�u ��H�� ]�@UH�� H��H�MP��N��H�� ]�@UH�� H��H�M@�E ��H�� ]�@UH�� H��H�MP��N��H�� ]�@UH�� H��H�M@� ��H�� ]�@UH�� H��H�M(�N��H�� ]�@UH�� H��H�Mp�����H�� ]�@UH�� H��H�MP�mN��H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��H�MP�HM��H�� ]�@UH�� H��H�M8�0M��H�� ]�@UH�� H��H�Mx�M��H�� ]�@UH�� H��H�M`� M��H�� ]�@UH�� H��H�Mx�=���H�� ]�@UH�� H��H�MP�%���H�� ]�@UH�� H��H�M0�L��H�� ]�@UH�� H��H�M0�����H�� ]�@UH�� H��H�M8�}M��H�� ]�@UH�� H��H�MP�����H�� ]�@UH�� H��H�M`����H�� ]�@UH�� H��H�Mx����H�� ]�@UH�� H��H�Mp�M��H�� ]�@UH�� H��H�Mp�M��H�� ]�@UH�� H��H�M@��L��H�� ]�@UH�� H��H�MP��L��H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��H�MP�L��H�� ]�@UH�� H��H�M@�����H�� ]�@UH�� H��H�M@���H�� ]�@UH�� H��H�M0�-���H�� ]�@UH�� H��E ����t�e �H�Mh����H�� ]�@UH�� H��H�M@�*K��H�� ]�@UH�� H��H�M@�K��H�� ]�@UH�� H��H�MH��J��H�� ]�@UH�� H��H�MH��J��H�� ]�@UH�� H��H�M@��J��H�� ]�@UH�� H��E ����t�e �H�Mp�J��H�� ]�@UH�� H��H�M@�J��H�� ]�@UH�� H��H�MX�tJ��H�� ]�@UH�� H��H�Mx�\J��H�� ]�@UH�� H��E(����t�e(�H���   �3J��H�� ]�@UH�� H��H��(  �J��H�� ]�@UH�� H��H���   ��I��H�� ]�@UH�� H��H���   ��I��H�� ]�@UH�� H��H���   ��I��H�� ]�@UH�� H��H��@  �J��H�� ]�@UH�� H��H��  �I��H�� ]�@UH�� H��H�MH�yI��H�� ]�@UH�� H��H���   �^I��H�� ]�@UH�� H��H���   �CI��H�� ]�@UH�� H��H���   �(I��H�� ]�@UH�� H��H�MP�J��H�� ]�@UH�� H��H�Mx��I��H�� ]�@UH�� H��H�M8��I��H�� ]�@UH�� H��H�M@�I��H�� ]�@UH�� H��H�MP�H��H�� ]�@UH�� H��H�Mp�H��H�� ]�@UH�� H��H���   �}H��H�� ]�@UH�� H��H�M8�eH��H�� ]�����@UH�� H��H�M`H������H�� ]�@UH�� H��H�M8����H�� ]�������������@UH�� H��H�M0�	H��H�� ]�@UH�� H��E ����t�e �H�M`��G��H�� ]���@UH�� H��H�MH��G��H�� ]���������@UH�� H��H�M@�H��H�� ]�@UH�� H��E ����t�e �H�Mx�xH��H�� ]���@UH�� H��H�M@辅��H�� ]�@UH�� H��E ����t�e �H���   蕅��H�� ]����������������@UH�� H��H�M8�H��H�� ]���������@UH�� H��H���   �;��H�� ]�@UH�� H��H�M0�#��H�� ]�@UH�� H��H�Mp���H�� ]������@UH�� H��E ����t�e �H�Mx� *��H�� ]�@UH�� H��H�MH�*��H�� ]�@UH�� H��E ����t�e �H�Mp��)��H�� ]�@UH�� H��H�MH��)��H�� ]�@UH�� H��E ����t�e �H���   �)��H�� ]�@UH�� H��H�MX�)��H�� ]�@UH�� H��E ����t�e �H�Mp��E��H�� ]�@UH�� H��H�MH��E��H�� ]������@UH�� H��H���   �����H�� ]������@UH�� H��H�M0�E��H�� ]�@UH�� H��E ����t�e �H�M`�cE��H�� ]�@UH�� H��H�MP�KE��H�� ]�@UH�� H��H�M8�3E��H�� ]�@UH�� H��H�M@�E��H�� ]�@UH�� H��E ����t�e �H�Mp��D��H�� ]�@UH�� H��H�M@��D��H�� ]�@UH�� H��E ����t�e �H�Mp�D��H�� ]�@UH�� H��H�M0����H�� ]�@UH�� H��E ����t�e �H�Mp�΂��H�� ]�@UH�� H��H�M0�VE��H�� ]�@UH�� H��E ����t�e �H�M`�0E��H�� ]�@UH�� H��H�M@�#D��H�� ]�@UH�� H��E ����t�e �H�Mp��C��H�� ]�@UH�� H��H�M@��C��H�� ]�@UH�� H��E ����t�e �H�Mp�C��H�� ]�@UH�� H��H�M@�����H�� ]�@UH�� H��E ����t�e �H���   �~C��H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��E ����t�e �H�M`����H�� ]�@UH�� H��H�MP�D��H�� ]�@UH�� H��H�M@�e���H�� ]�@UH�� H��E ����t�e �H���   ��C��H�� ]�@UH�� H��H�MP��B��H�� ]�@UH�� H��E0����t�e0�H���   �B��H�� ]�@UH�� H��H�MP�����H�� ]�@UH�� H��E0����t�e0�H�Mp����H�� ]�@UH�� H��H�M8�EC��H�� ]�@UH�� H��E ����t�e �H���   �'B��H�� ]�@UH�� H��H�MP�C��H�� ]�@UH�� H��H�M@�L���H�� ]�@UH�� H��E ����t�e �H���   ��A��H�� ]�@UH�� H��H�MP�B��H�� ]�@UH�� H��H�M@�����H�� ]�@UH�� H��H�MP�{B��H�� ]�@UH�� H��H�M@�����H�� ]�@UH�� H��H�MP�KB��H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��H�M@�B��H�� ]�@UH�� H��E ����t�e �H�Mp��A��H�� ]����������������@UH�� H��H�M@��A��H�� ]�@UH�� H��E ����t�e �H�Mx�A��H�� ]�@UH�� H��H�M@�A��H�� ]�@UH�� H��E ����t�e �H�Mx�jA��H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H�MX��#��H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H�M8�#��H�� ]�@UH�� H��H�MH�R���H�� ]�@UH�� H��H�MX�j#��H�� ]�@UH�� H��E$����t�e$�H���   �~��H�� ]�@UH�� H��H�MH�����H�� ]�@UH�� H��H�MX�#��H�� ]�@UH�� H��E$����t�e$�H���   �}��H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H�M8�"��H�� ]�@UH�� H��H�MH�p���H�� ]�@UH�� H��H�M8�"��H�� ]�@UH�� H��H�MP�@���H�� ]�@UH�� H��H�M`�X"��H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H�M8�("��H�� ]�@UH�� H��H�MH�����H�� ]�@UH�� H��H�MX��!��H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H�M8��!��H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��H�MP�!��H�� ]�@UH�� H��H�MH�P���H�� ]�@UH�� H��H�M8�h!��H�� ]�@UH�� H��H�M@� ���H�� ]�@UH�� H��H�MP�8!��H�� ]�@UH�� H��H�MH�����H�� ]�@UH�� H��H�M8�!��H�� ]�@UH�� H��H�M@�����H�� ]�@UH�� H��H�MP�� ��H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H�M8� ��H�� ]�@UH�� H��H�M@�`���H�� ]�@UH�� H��H�MP�x ��H�� ]�@UH�� H��H�MH�0���H�� ]�@UH�� H��H�M8�H ��H�� ]�@UH�� H��H�MH� ���H�� ]�@UH�� H��H�MX� ��H�� ]�@UH�� H��H�MH�����H�� ]�@UH�� H��H�M8����H�� ]�@UH�� H��H�M@����H�� ]�@UH�� H��H�MP���H�� ]�@UH�� H��H�MH�p���H�� ]�@UH�� H��H�M8���H�� ]�@UH�� H��H�MH�@���H�� ]�@UH�� H��H�MX�X��H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H�M8�(��H�� ]�@UH�� H��H�MH�����H�� ]�@UH�� H��H�MX����H�� ]�@UH�� H��H�MH����H�� ]�@UH�� H��H�M8����H�� ]�@UH�� H��H���   �<��H�� ]�@UH�� H��H�MP��?��H�� ]�@UH�� H��H�M8�?��H�� ]�@UH�� H��H�M(�ծ��H�� ]�@UH�� H��H�M8�}?��H�� ]�@UH�� H��H�M(襮��H�� ]����������������@UH�� H��H�M@�����H�� ]�@UH�� H��H�MP����H�� ]�@UH�� H��E ����t�e �H�Mx����H�� ]�����������@UH�� H��H���   �&:��H�� ]�@UH�� H��H��   �:��H�� ]�@UH�� H��E0����t�e0�H���  ��9��H�� ]�@UH�� H��H���   ��9��H�� ]�@UH�� H��H��P  �9��H�� ]�@UH�� H��H��  �9��H�� ]�@UH�� H��H���   �v9��H�� ]�@UH�� H��H��h  �[9��H�� ]�@UH�� H��H��8  �@9��H�� ]�@UH�� H��H�M8�(9��H�� ]�@UH�� H��H�M8�9��H�� ]����������������@UH�� H��H�MP��8��H�� ]�@UH�� H��E0����t�e0�H���   ��8��H�� ]����������������@UH�� H��H�M(H�E(H� � �E$H�E(�M$H�������H�� ]��@UH�� H���]	 ����H�� ]��������@UH�� H��   �O���H�� ]�������@UH�� H��}  uL�MXD�EPH�UHH�M@����H�� ]������@UH�� H��H�M H�E H������H�� ]�����������������@UH�� H��H�MHH�EHH� � �E(�E(=  �u	�E$   ��E$    �E$H�� ]�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@WH��H�$H��3��   �H��_���������������������@WH��H�$H��3��   �H��_���������������������H��(H�-�  ��@��H�9  �����H��(����������������@WH��H�$H��3��   �H��_�����@WH��H�$H��3��   �H��_�����@WH��H�$H��3��   �H��_�����@WH��H�$H��3��   �H��_�����@WH��H�$H��3��   �H��_�����@WH��H�$H��3��   �H��_�����H��(3�H�c�  ����H��(����������@WH��H�$H��3��   �H��_�����H��(�W����e�  H��(�������������H��(�   �   ������   ��������    ��������  H��(�����������@WH��H�$H��3��   �H��_�����@WH��H�$H��3��   �H��_�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������H��(H���  ��.��H��(����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ���           ���            ��   0��   P��   p��   ���   ���   ���   ���   ��   ���   P��   0��   ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           0��                                                                                                                                                                                                                                                                           P��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               i{�Q       s   t\ tF     i{�Q          �\ �F                �������N���������������C-DT�!	@-DT�!�?                                       Ocontainer.png  Ocontainer  �������N    ���������������C-DT�!	@-DT�!�?"�   �k            l `                                  "�   �j            �j 8                  "�   tl            |l 8                  "�   �l            �l �                  "�   xm            �m H                  ^�   
 �   �� �    � �    � �   @� �   `� �   �� �   �� �   �� �   �� �    � �    � �   @� �   `� �   �� �   �� �   �� �                                    _�    �   �� �    � �    � �   @� �   `� �   �� �   �� �   �� �   �� �    � �    � �   @� �   `� �   �� �   �� �   �� �   ���   ���   ��   0��   ���    ��    ��   @��   `��   ���   ���   ���   ���    ��    ��   @��                                                                   �_�   i �   # �   � �   A �   s �   � �   x �   �� �   �� �   �� �    � �    � �   @� �   `� �   �� �   �� �   �� �   ���   ���   ��   0��   ���    ��    ��   @��   `��   ���   ���   ���   ���    ��    ��   @��                                                           src/ContainerObject.cpp         333333�?        ffffff�?              �?             �o@        ../../resource/_api/c4d_resource.cpp    ../../resource/_api/c4d_resource.cpp    #   #   #   #   #   #   #   #   #   #   M_EDITOR        M_EDITOR        "�   �n            �n 8          "�   �n            �n @          "�   @o            Xo X          "�   �o            �o x          "�   `p            �p �          "�   8q            hq �          "�   Xr            pr �          "�   �r            �r �          "�   hs            xs 8          "�   �s            �s 8          H`�   �L �   �������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_file.cpp        ../../resource/_api/c4d_file.cpp        "�   �t            �t            "�   �t            �t            "�    u            (u            "�   Xu            `u            "�   �u            �u            "�   �u            �u 8          "�   0v            @v 8          "�   xv            �v 8          "�   �v            �v 8          "�   `w            pw (          "�   �w            �w 8          "�   �x            �x (          "�    y            y @          "�   �y            �y 8          "�   �z            �z 8          "�   �z            �z 8          "�   0{            @{ 8          "�    ~         	   (~ 0          "�   �~            �~ 8          "�                 8          "�   P            h X          "�   �            � 8          "�    �            0� 8          res �������N    ���������������C-DT�!	@-DT�!�?"�   p�            �� h          ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  �������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  "�   ��            � 8          "�   ��            Ȅ 8          "�   ��            �� 8          "�   0�            8�            "�   h�            p�            "�   ��            �� 8          "�   h�            x� @                          p:\applications\maxon\cinema 4d r14.041\resource\_api\c4d_misc/datastructures/basearray.h       Progress Thread 0%      ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp %   ����../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ���N~   ���������������C-DT�!	@-DT�!�?"�   H�            P� @          "�   ؊            �� 0          "�   ��            �� X          "�   P�            `� 8          "�   ��            �� 8          "�   �            (� h          "�   p�            �� 8          "�   Ѝ            ؍ H          "�   D�            L� 0          "�   ̎            ܎ X          "�   $�            4� H          "�   ��            �� (          "�   �            � (          "�   d�         	   �� p          "�   ��            �� h          "�   ��            �� h          "�   ܓ            � 8          "�   �            ,� 8          "�   t�            �� 8          "�   4�            <�            "�   t�            �� (          "�   ܕ            � 8          "�   �            � 8          "�   \�            d� @          "�   ��            �� @          "�   �            �� 8          "�   4�            T� p          "�   ܗ            � �          "�   ��            �� 0          "�   �         	   � x          "�   ��            �� P          "�   ��            �� X          "�   \�            t� h          "�   Ԛ            ܚ `          "�   ��            �� (          "�   ܛ            � 8          "�   0�            @� 8          "�   ��            �� 0          "�    �            (�            ha�   �h�   �� �   �� �    � �    � �   @� �   �� �   �� �   � �   0� �   P� �   @a�   ph�    � �   @� �   `� �   �� �   �� �   �� �   �� �   �� �   �a�   �h�    � �   @� �   `� �   �� �   �� �   �� �   �� �   P>�   p`�   pi�    � �   @� �   `� �   �� �   �� �   �� �   �� �   �D�   `b�   �i�    � �   @� �   `� �   �� �   �� �   �� �   �� �    F�   pF�   �F�   �F�   �F�   �F�   �F�   �F�   �F�   PG�   �G�   �G�   H�           -DT�!	@      Y@     �f@     @�@�������������        ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  nncnt<ncnt  ����../../resource/_api/c4d_baseobject.cpp  %s(%d): %s  ���N../../resource/_api/c4d_baseobject.cpp  nncnt==ncnt     ../../resource/_api/c4d_baseobject.cpp  %s(%d): %s      ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ���������������C-DT�!	@-DT�!�?"�   p�            x� 0          �b�   P��   ���           p:\applications\maxon\cinema 4d r14.041\resource\_api\c4d_misc/datastructures/sort.h    Stop:   Stop    ����MbP?�������N���������������C-DT�!	@-DT�!�?"�   $�            ,� @          "�   l�            t� (          "�   ��            �� H          �������?-DT�!�?      �-DT�!��       �       �"�   �            � @          "�   ��            �� @          "�   ��            �� @          "�   T�            d� @          "�   Ĩ            ̨ `          ../../resource/_api/c4d_pmain.cpp       ../../resource/_api/c4d_pmain.cpp       %s     "�   Ī            Ԫ (          "�   \�            t� 0          "�   ī            ԫ 8          "�   �            � 8          "�   �            �� (          "�   \�            l� (          "�   8�            H� 8          "�   ��            �� 8          "�   0�            @� 8          "�    �            � 8          "�   H�            h� 8          "�   ذ            � H          "�    �            0� H          "�   h�            p�            "�   ��            �� 8          "�   �            0� 8          "�   ��            �� 8          "�   �            �� 8          "�   г            � 8                  p:\applications\maxon\cinema 4d r14.041\resource\_api\c4d_general.h     ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp          �?   ����A  4&�kC �Ngm��C  4&�k�`c�   �R�    S�   ���   ���   �������N���������������C-DT�!	@-DT�!�?"�    �            0� 8          "�   h�            x� 8          "�   ��            �� 0          "�   �            (�            "�   p�            �� 0          "�   �             � 0          "�   `�            p�            "�   ��            ȹ            "�   �             � 8          "�   x�            ��            "�   к            � 0          "�   8�            H�            "�   ��            �� (          "�   ��            �            "�   X�            h� (          "�   ��            м            "�   4�            D� (          "�   ��            ��            "�   ��            � (          "�   `�            p�            "�   ��            Ⱦ 0          "�    �            0�            "�   |�            �� (          "�   �            ��            "�   <�            L� 0          "�   ��            ��            "�   ��            � 0          "�   d�            t�            "�   ��            � �          "�   ��            �� 0          "�   ��            � 0          %H:%M:%S         [%s %s L%d]    WARNING:    
   CRITICAL:   �������N    ���������������C-DT�!	@-DT�!�?%s      ../../resource/_api/c4d_misc/memory/debugglobals.cpp    ../../resource/_api/c4d_libs/lib_ngon.cpp       ../../resource/_api/c4d_libs/lib_ngon.cpp       ../../resource/_api/c4d_libs/lib_ngon.cpp       ../../resource/_api/c4d_libs/lib_ngon.cpp       ../../resource/_api/c4d_libs/lib_ngon.cpp       ../../resource/_api/c4d_libs/lib_ngon.cpp       ../../resource/_api/c4d_libs/lib_ngon.cpp       "�   �            0� (          no baselist  GB  MB  KB  B      ../../resource/_api/c4d_string.cpp      "�	   ��            �� �          "�   ��             � 0          "�   0�            8� 0          "�   @�            P� H                �@�c�   ���           f:\dd\vctools\crt_bld\self_64_amd64\crt\src\crtdll.c    ( _ _ o n e x i t e n d   ! =   N U L L   & &   _ _ o n e x i t e n d   ! =   N U L L )   | |   ( _ _ o n e x i t e n d   = =   N U L L   & &   _ _ o n e x i t e n d   = =   N U L L )     % s                 f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ 6 4 _ a m d 6 4 \ c r t \ s r c \ a t o n e x i t . c     f:\dd\vctools\crt_bld\self_64_amd64\crt\src\atonexit.c  ���   @��                       p                                                                                       ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       RSDS#ိ��zA�z&���`   P:\applications\MAXON\CINEMA 4D R14.041\plugins\c4dpl-container-object\containerobject.pdb      -   -                                                                                                                                                                                                                                                                                                                   � H^ ^                                    `^         x^ �^                  �        ����    @   H^                     (�         ����    @   �^                                �^         �^                        P� 0_  _                                    H_         p_ x^ �^                             P�        ����    @   0_                                x� �_ �_                                    �_         ` p_ x^ �^                                 x�        ����    @   �_                                (� �^ H`                            �� �` p`                            �`         �` �`                 ��        ����    @   �`             ��         ����    @   a                        0a         �`                        �� a @a                            �� �a ha                            �a         �a             ��         ����    @   �a                        � b �a                             b         8b �`                 �        ����    @   b                        8� �b `b                            �b         �b �` �`                     8�        ����    @   �b                        `� c �b                            (c         8c             `�         ����    @   c                        �� �c `c                            �c         �c             ��         ����    @   �c                        ��  d �c                            d         (d             ��         ����    @    d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      B  	 	B  	 	B   B   b       p	 	B   B   B  	 	B   �  b�  )     ����8�      �     �  ����D     ^           2P 2P B   B   B   �p`       B   B   B  	 	B  	 	B  	 	B  	 	B  	 	B   B   p	 	B  	 	B   b   b  	 	B  	 	B  	 	B   B   �   b    b� �( ������     �� ������    �� �  �����      �     '     w     �  ���� 2P 2P 2P                 �  b� P)     ����� }  �����      �  ����     2P" # b� �)     ����p�     ��     �� ������     �  �����       �   ����"      2"     E"      n"     �"      �#  ����C$     W$  ����l$                   2P 2P 2P 2P  b� �)     ���� � �����     �  ����z+      �+  �����+     �+  ����     2P 2P   �   B   b   �   b   �  	 	B  	 	B   B   b  	 	b  	 	B   B  	 	B   B   B   B   b   b   B   B   B   b   B  	 	B   	�  b�  . ����@� p3  �����3      �3  ���� 2P �  b� H. ����X� �3  ����4      G4  ���� 2P	 	b   B  	 	B  	 	�   B    b� p. ������     ��    �� �6  ����77     L7     �7     �7      �7     8       2P 2P 2P#  b� �. �����     ݸ    ��    6� @8  �����8     �8     �8     9      9     i9     �9     �9      �9     9:       2P 2P 2P 2P&  b� �. ������     Q�    i�    ��    ¹ `:  �����:     �:     �:     %;      <;     �;     �;     �;      <     Q<     �<     �<      �<     !=       2P 2P 2P 2P 2P&  b� �. �����     ݹ    ��    6�    Q�    l� P=  �����=     �=     �=     >      ,>     |>     �>     �>      �>     J?     �?     �?      �?     @     Q@     @      �@     �@       2P 2P 2P 2P 2P 2P b  	 	B   �    b� / ������ ������    ˺ `B  �����B      �B  ����IC     �C     �C     �C  ���� 2P 2P 2P  b� 8/ ������ �����    8� 0D  �����D      �D  ����2E     iE     �E     �E  ���� 2P 2P 2P B   B  	 	B  	 	B  ! �  b� `/ ������     p� H  ����sH     �H       2P 2P B   B  	 	�  	 	B  	 	B   �  b� �/ ����Ȼ     �� @J  �����J     �J       2P 2P	 	B   B  	 	B   B   B   B  	 	B   B   B   B   B   B   B   B   B   B  	 	B   B   	b  b� 80 ���� � �M  �����M      �M  ���� 2P b  b� `0 ����� �M  ����N      GN  ���� 2P b  b� �0 ����0� `N  �����N      �N  ���� 2P b  b� �0 ����H� �N  �����N      'O  ���� 2P 	b  b� �0 ����`� @O  ����RO      iO  ���� 2P B   b  	 	B   �  b�  1 ������     x� PP  �����P     �P       2P 2P B   �  b� (1 ����μ     �� Q  ����YQ     vQ       2P 2P �  b� P1 �����     �� �Q  �����Q     R       2P 2P �  b� x1 ����P�     8� 0R  ����pR     �R       2P 2P	 	B  	 	B   B   B   B   B   B   B   B  	 	B   B   �  b� �1 ������     y� @U  ����tU     �U       2P 2P B   B   b   �  b� �1 ����Ͻ     �� �V  �����V     W       2P 2P �  	 	B   B   B   B   B   B  	 	B  	 	B  	 	B   B   B   B   B   B   B   B   B   B   B   B   �  b� �1 ������ @\  ����b\      }\  �����\      �\  ���� 2P b   �  b� 2 �����  ]  �����]      �]  ���� 2P b   b   b   b   B   B   B   B   B   B   B   B   B   B   �  b� @2 ����%� �b  ����%c      8c  ���� 2P b   �   b   b   b   b   B  	 	B   �   b   B  	 	B   B  	 	B  	 	B  	 	B  	 	B  	 	B  	 	B   B   �  b� h2 ����U�     =� j  ����Yj     vj       2P 2P B  	 	B  	 	B  	 	B   �  b� �2 ������     ~� `k  �����k     �k       2P 2P �  b� �2 ����׾     �� �k  ����Fl     `l       2P 2P B  	 	B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   b   B   B   B   B   b   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   B   b   B   b  	 	B   B   B   B   B  	 	B   B  	 	B  	 	B  	 	B  	 	B   B  	 	B   b  	 	B   b   B   B   B   B   B   B   B  	 	B   	�  b� �2 ������ 0�  ����R�      h�  ����{�      ��  ������      ݁  �����      ��  ���� 2P	 	B   B   b   B  	 	B   B   	�  b� 3 ����-�     � ��  ����܃     ��       2P 2P 	�  b� 03 ����n�     V�  �  ����_�     |�       2P 2P	 	b    b� X3 �����     ��    �� ��  ����*�     A�  ����Z�     ��     ��       2P 2P 2P �  b� �3 ����'�     � ��  ����:�     W�       2P 2P B   B  	 	B   �  b� �3 ����h�     P� 0�  ������     ��       2P 2P B   B   p B   B   B   B   B   B   B   B  	 	B   b   B   B  	 	B   B   B  	 	B   B   B  	 	B   b   �   b  	 	B   B  	 	B   B   B  	 	B   B   B   B   B  	 	B  	 	B   B  	 	B   B  	 	B  	 	B   B   b   B   B   B   B   B  	 	B   B   B   B   B   B  	 	B   B  	 	B   B   b   B   b   B   B   /  + b�  4 ������     ��    ��    ��    ��    � @�  ������      ��     ɞ     �     �     7�     u�     ��     ��     ��     ��      ��  ���� 2P 2P 2P 2P 2P 2P B  	 	B   B   p B  	 	B  	 	B  	 	b  	 	B   p "   b   B  	 	B   B   B   b   b   B   B   B   B   �  b� h5 ����H�     0� ��  ������     �       2P 2P	 	B  	 	B   B   B   B   B   B   B   B  	 	B   b   b  	 	B   b   B  	 	B   	�  b� �5 ����n� ��  �����      �  ���� 2P b   B   b   b   b   b   �   �   �   B   B  	 	B  	 	B  	 	B   B   B  	 	B   B  ! �  b� �5 ������     �� ��  �����     �       2P 2P B  	 	B   b  	 	B   b   �   B  	 	B  	 	B   B   B  	 	B   	b  b� �5 ������ `�  ������      ��  ���� 2P 	b  b� 6 ������ ��  ������      ��  ���� 2P	 	b   �  b� 06 ������ �  �����      <�  ���� 2P	 	�   �  	 	B   b   �   B  	 	B   B   B  	 	B   b   b  	 	b   b   �   b   b    b� X6 ����(� ����@�  �  ����U�      ��  ������     ӽ  ���� 2P 2P b   b   �   �   b   b   �   B   B  	 	"   b   �  	 	"   b   �   b   B   b  	 	b   B   b  	 	b  
 
B   "   b  	 	B   �  b� h= ������     �� �g �����g    �g      2P 2P b   b   B   B  	 	B  	 	B   B  	 	B  	 	B  	 	B  	 	B   b   b   �    b� 8 ����`� ��  ������      ��  ���� 2P B  	 	B  	 	B  	 	B  	 	B  	 	B   B   B   B  	 	B   B   B   B   B   B   B   B   B   �   b   B   B   b   b   �   b   �   �   B   B   B  	 	B  	 	B   B   b  	 	B  	 	B   b   �   B   B   B   B   	�  b� @8 ����x� @�  ����p�      ��  ���� 2P B   B   b   B   b   b   �   b   B  	 	B  	 	B  	 	B  	 	B   b   �  	 	B   B  ! �  b� h8 ������     �� @�  ������      ��  �����     ,�       2P 2P B  	 	b  	 	�  	 	�   B   �   B   B  	 	B   b   b   �  ! �  b� �8 ������     �� ��  ������      ��     ��      ��  ���� 2P 2P# �  b� �8 �����     �  �  ����S�      ��     ��      ��  ���� 2P 2P �   �   �  $  b� �8 ����1�     I�  �  ������      +�     9�      D�  ���� 2P 2P! �  b� 9 ����a�     y� `�  ������      �     �      �  ���� 2P 2P �  ! �  b� 09 ������ ��  ����"�      P�  ���� 2P �   b   b   B   �   �   �p`   �  b� X9 ������  �  ����'�      N�  ����^�      u�  ���� 2P �   B   �   �   �   �   �   �  $  b� �9 ������     �� � �����     +    W     b ���� 2P 2P$  b� �9 ������     	� � �����     �          ���� 2P 2P �   b   b   b   �   �  ! �  b� �9 ����!� 0 ����\     � ���� 2P! �  b� �9 ����9� � �����      ���� 2P �   b   �   �   �   �   �   �   �  $  b�  : ����Q�     i�     ��     �� � ����     &    ;     W    l     �    �     � ���� 2P 2P 2P 2P b  	 	�   B   B   B   B   �   �   �   b   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   b   �   �   �   �   b   �  	 	�   B   �  	 	B   B   b   B   b    b� H: ������ �( ����
)     �) ���� 2P �   �   B   B   b   b   b   �   �   �   �   �   �   �   �  	 	�   �  	 	�   �   �  	 	�  	 	�   �  	 	�   b  #  b� p: ������ �6 �����6     ]7 ���� 2P	 	b   �   �   b   �  b� �: ������ `: �����:     �: ���� 2P	 	B   �  b� �: ������     � p; �����;     �;    �;     �; ���� 2P 2P �  b� �: ����)�     A�  < ����g<     �<    �<     �< ���� 2P 2P	 	B  	 	B   �   B   b   �   �   �   �   �  	 	B  	 	B   b   b  b� ; ����Y� PE ����wE     �E ���� 2P b   �  b� 8; ������     q� �F ����G    4G      2P 2P	 	"   B  	 	B   b   �  b� `; ������ �H �����H     �H ���� 2P �  b� �; ������ I ����eI     vI ���� 2P	 	b   b   �  b� �; ������ @J �����J     �J ���� 2P �  b� �; ������ �J ����8K     gK ���� 2P B   B   b  	 	B   �  b�  < ����'�     � �L �����L    �L      2P 2P  b� (< ������     M�    e�    }�  M ����MM    �M    �M    	N    N    EN      2P 2P 2P 2P B   b   B  	 	B   - b� P< ������ ������ ������ ����� ����*�    E� �O ����P     $P ����PP    �P �����P    -Q ����lQ    �Q �����Q    +R    nR    |R ���� 2P 2P 2P 2P 2P 2P 	�  b� x< ����`� �R ����pS     �S ���� 2P  b� �< ����x�     ��    �� ������ �S ����T     HT    qT    �T    �T     �T �����T    �U ���� 2P 2P 2P 2P  b� �< ������ ������  V ����uV     �V ����W    fW ���� 2P 2P b  	 	B   b   �  b� �< ����� 0Z ����_Z     �Z �����Z     �Z �����Z     P[ ���� 2P b   �    b� = ����)�     A�    Y� p\ �����\     �\    �\    �\    ]     @] ���� 2P 2P 2P$  b� @= ����t� `] �����]     ^ ����^     T^ ���� 2P b   �   b   �    p`  p` �p`   �p`   B   B   B   B  	 	B   B   B  	 	B   B   B   B   B   B   B  ! �  b� �= ������     p� @n �����n    �n      2P 2P bp`   �  b� �= ����H�     0� @m �����m    �m      2P 2P B   B   B   B   B   	�  b� �= ������     ��  d ����$d     Hd    _d     jd ���� 2P 2P	 	B   B   p	 	"  	 	"   b  b� > ����� l ����'l     �l ���� 2P	 	"  	 	"   Bp`  	 	"   Bp`  	 	B   B   B   B  	 	B  	 	B   B  	 	B   B  	 	B   B  	 	B   B  	 	b   B  	 	B   B   B   B   B   B  	 	B   b   b   B   B   B  	 	B   b  ! �  b� �B ������ �y ����Oz     �z ���� 2P	 	B   B   B  	 	B   B  	 	B   �   b  	 	B  	 	B   B  	 	B  	 	B  	 	B  	 	B  	 	B   �p`  	 	B   B   B   B   B   B   b   �   B  	 	B  	 	B  	 	B   B   B   B   B   B   b  	 	B  	 	B  	 	B  	 	B  	 	B  	 	B   B   B   b   b   �   �  	 	B   B   B  	 	B  	 	B   B   B  	 	B   B  	 	B   B   B   B   B   B   B  	 	B   b  	 	B   B   B  	 	B   B   B  	 	B  	 	b  	 	B   �p`   �p`  	 	B   B   B   B  	 	B   b   b  	 	B   b  	 	B   B   1 p` B   B   �   �   B   B   �  	 	B   b  	 	B   �   �   b   B     b   B  	 	B   �   �  	 	B   B  	 	B   B   B   B   B   B   B   B   B  	 	B  	 	B  	 	B  	 	B  	 	B  	 	B  	 	B   b   B   B   B   p b  	 	"   B   B  	 	b   "   "   B   B   B   �   B  ' �  P� `   ' �  P� @   ' b  P� (   " �  P� 0    B   �   b  
 
B  
 
B  
 
B   b  	 	B   b   b   b   b    p` B    p` b   b    p` �p`   � p`$ ! b� hC ������ �� ����x�     �� ������     �� ���� 2P$ # b� �C ������ 0� ������     � �����     y� ���� 2P& 7 p`b� �C ����� �� ���� �     �� ���� 2P O  b  	 	b   B   p	 	B    p`  p` B  	 	B   �p`   �p`   �p`   B   B   B   B   "   b  	 	b   b   �   b   b   b  	 	b   b   b  	 	b   b   b   b   b   �  b� D ����0�     V� p� ������     �� ����
�    $�      2P 2P b   b  	 	b   b   �   �  b� 8D ����n�     �� �� ������     �� ����(�    B�      2P 2P b  	 	b   b   b   b  	 	b  	 	b   b   b   b  	 	b   �   b   b   b   b   b  	 	b   b   b   b   b   �  	 	b   b   �  b� `D ������     �� @ �����     � �����          2P 2P b   b   b   b  	 	b   b   b   b  	 	b   b   �  b� �D ������     � 	 ����Q	     c	 �����	    �	      2P 2P B   B   �  #  b� �D ����0� �
 �����
      ����!     � ���� 2P b   b   B   b   b   B  	 	B   B   B   B   �   "  	 	B   B  	 	B   B   B  	 	B   B   B   b   B   B   b   b   b   B   B  	 	B   B   B  	 	B   B   B  	 	B   �   b   B  	 	B   B   B  	 	B   B   b   B   B   B   B   B   B   �   B   B   B   �   	�  b� 0E ����h�     P�  ����5    b      2P 2P B   B   B   B   B   B  	 	B  	 	B   b  	 	B   	�  b� XE ������     �� ������ � �����     �    � ���� 2P 2P B  	 	B   	�  b� �E ������     �� � �����    �      2P 2P 	�  b� �E �����     ��    ����?     Y       2P 2P B   B   B   B   B   B  	 	B  	 	B   B   B   B   B   B  	 	B   B   B   B   B   B   �  b� �E ����R�     :� `$ �����$    �$      2P 2P B   B   B   B   B   	�  b� �E ������     x� & ����5&    e&      2P 2P B  	 	B   �p
`   B   B   B   B   B   B   B   B   B   B   B   b   B  	 	B  	 	B   �  b�  F ������     �� �* ����+    !+      2P 2P �  b� HF �����     �� @+ �����+    �+      2P 2P	 	B  	 	B  	 	b  	 	b  	 	b   B   B   B   B   B  	 	B   B   B   �  b� pF ����J�     2� �. �����.    /      2P 2P	 	B   B   B   B  - 	P� 0  	 	b   �   �   �  	 	B   B   b  	 	B   b   B  	 	B    �  b� �F ������     s� �4 �����4    5      2P 2P 	�  b� �F ������     ��    ��     ��  5 ����X5    p5    �5     �5    �5      2P 2P 2P	 	B   �   �  ! �  b� �F ����"�     
�  7 �����7    �7      2P 2P! �  b� G ����c�     K� �7 ����P8    j8      2P 2P �  b� 8G ������ �8 �����8     
9 ���� 2P �  b� `G ������     ��    ��  9 ����U9     m9 ����}9    �9    �9    �9      2P 2P 2P �  b� �G ������     #�    ;� : ����E:     ]: ����m:    �:    �:    �:      2P 2P 2P �  b� �G ����S�     k�  ; ����.;     k;    y;     �; ���� 2P 2P �  b� �G ������     �� �; �����;     <    <     $< ���� 2P 2P b   b   B  	 	B  	 	B  	 	B   B   B   B   B   B   �   B   B   B   B   B   B   �  b�  H ������     �� �@ �����@    A      2P 2P	 	B   B   B  	 	B   B   B   B   B  	 	B   B  	 	B  	 	B   B   B   �   B  	 	B  	 	B   b   B  
 
B  	 	�   B   b   B   b  	 	B  	 	B  	 	B  	 	B   B   B   B  	 	B   �   B   b  	 	B  	 	B  	 	B   B  	 	B   B  	 	B  	 	B   B   B   B  	 	B  	 	B  	 	B   B   B   B   B  	 	B  	 	B   B   b  	 	B   B   B  	 	B   B  	 	B   �  b� hI �����      � `U �����U    �U      2P 2P B   B  	 	B  	 	B  	 	B   B   B   B   b  	 	B  	 	B  	 	B  	 	B   B   B   B   b   B   B   B   B   B   B   B   B  	 	B   B   B   B   B   B  	 	B   �  b� �I ����V�     >�  ^ ����y^    �^      2P 2P 	�  b� �I ����|�     �� �^ �����^     �^    #_     >_ ����N_     \_ ���� 2P 2P 	�  b� �I ������     �� �_ �����_     �_    �_     �_ ���� 2P 2P �  b� J �����     ��    ��  ` ����*`    G`    �`    �`     �`    �`      2P 2P 2P �  b� 0J ����e�     5�    M� a ����:a    Wa    �a    �a     �a    �a      2P 2P 2P �  b� XJ ������     ��  b ����Gb     db    b     �b ���� 2P 2P �  b� �J ������     �� �b �����b     �b    �b     
c ���� 2P 2P 	�  b� �J ������     �  c ����=c     Zc    �c     �c �����c     �c ���� 2P 2P �  b� �J �����     6� �c ����d     6d    Qd     \d ���� 2P 2P 	�  b� �J ����N�     f� �d �����d     �d    �d     e ����e     ,e ���� 2P 2P �  b�  K ����~�     �� Pe ����ue     �e    �e     �e ���� 2P 2P �p`  b� HK ������     �� �e �����e     f    Jf     kf ����f     �f ���� 2P 2P �  b� pK ������     �� �f �����f     g    g     *g ���� 2P 2P �p`  b� �K �����     &� @g ����dg     �g    �g     �g �����g     h ���� 2P 2P �  b� �K ����>�     V� 0h ����Wh     th    �h     �h ���� 2P 2P bp`   bp`   �p`  b� �K ����n�     �� pi �����i     �i    �i     j ����j     ;j ���� 2P 2P �  b� L ������     �� `j �����j     �j    �j     �j ���� 2P 2P �p`  b� 8L ������     �� �j ����k     !k    Zk     {k �����k     �k ���� 2P 2P �  b� `L ������     � �k �����k     l    /l     :l ���� 2P 2P 	�  b� �L ����.�     F� Pl ����ml     �l    �l     �l �����l     �l ���� 2P 2P �  b� �L ����^�     v�  m ����Em     bm    }m     �m ���� 2P 2P �p`  b� �L ������     �� �m �����m     �m    n     ;n ����On     kn ���� 2P 2P �  b�  M ������     �� �n �����n     �n    �n     �n ���� 2P 2P 	�  b� (M ������     � o ����-o     Jo    �o     �o �����o     �o ���� 2P 2P �  b� PM �����     6� �o ����p     "p    =p     Hp ���� 2P 2P 	�  b� xM ����N�     f� `p ����}p     �p    �p     �p �����p     q ���� 2P 2P �  b� �M ����~�     �� 0q ����Uq     rq    �q     �q ���� 2P 2P	 	b  	 	B  	 	B   B   B   B  	 	B   B    b� �M ������     �� �s ����t     )t    Ju     Uu ����iu    �u     �u ���� 2P 2P	 	B  	 	B   B  	 	B  	 	B   B   B  	 	B  	 	B  	 	B   b   B   b   B   b  	 	B   B   B   B   B   B   B   B  	 	B   �   B   B  	 	B  	 	B  	 	B  	 	B   �   �   B   B   �   	�  b� �M ������     �� � �����     �    :�     E� ����U�    ��     �� ���� 2P 2P 	�  b� N �����     )� Ѐ �����     ��    �     %� ����5�    ��     �� ���� 2P 2P B   B   B   B  	 	B   B   B   b   p	 	B  	 	B  	 	B   B  	 	B  	 	B  	 	B  	 	B  	 	B   B  	 	B  	 	B  	 	B  	 	B  	 	B   B  	 	B  	 	B  	 	B  	 	B  	 	B  	 	B  	 	B  	 	B   B  	 	B  	 	B  	 	B   B  	 	B  	 	B  	 	B   B  	 	B   �p`   �p`   �p`    p` B   B   B   B   B   B   B  	 	B  	 	B  	 	B   B   B  	 	B  	 	b   B  	 	B   b   B  	 	B  	 	B  	 	B   B   B   B  	 	B   B   B   b   B   B   B   B  	 	B   B   B   �   �   B  	 	B   p, 	P� 0   b  	 	B  	 	B  # � P� �   B  	 	B   �   B   B   b   b  	 	B   B   B   B   b  	 	B   b   �   [ p` b   b     �  	 	b   b   b   b  	 	b  	 	b  	 	b   b  	 	b   b   b   b   b   b   b  	 	b  	 	b   b   b  	 	b   b   b   b   b  	 	b  	 	b  	 	b  	 	b  	 	b   b   b   �   b   b   b   b   b   b   �   �   �   b   b   b   b   B  	 	b   �p`   p`  p` B   B  	 	B   b   b   B   b   B   B   B   B   �p`   �p`   �  b� 8P ������     P�    h� p� ������    ��    ��    ��      2P 2P 2P b   B   B  	 	B   �   �     �   �   B   B   B   �   �   �   b   b   B   B   b   B   b   B   b  " �  b�  Q �����     �� �� ����-�    J�      2P 2P �   �  P� P    1 b� �P ������     ��    ��     �    *�     E�    `�     {�    �� @� ������    ��    �    )�     H� ������    ��    ��    �     +� ����l�    ��    ��    ��     � ����.�    Q�    s�    ��      2P 2P 2P 2P 2P 2P 2P 2P 2P	 	B  	 	B  	 	B   	�  b� �P ������ �� ������     �� ���� 2P 	�  b� �P ������ � ����@�     [� ���� 2P B   p B     b   b  ��    �� � @� � �� � p�      2P 2P B  	 	b  	 	�  ��    ~� �� ��      2P �   �   B      B   b   B  	 	B  	 	b   b  ��    Q� �� ��      2P	 b  ��    � ;� �� ;�  2P	 	b  	 	B   B  		 	�  ��    %� �� � ��  2P �  
 
4 
2p
 
4 
2p B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  i{�Q    �          � � � � &�   containerobject.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  XQ�           .?AVNodeData@@          XQ�           .?AVBaseData@@          XQ�           .?AVObjectData@@        XQ�           .?AVContainerObject@@           XQ�           .?AVSubDialog@@ XQ�           .?AVGeDialog@@  XQ�           .?AVGeUserArea@@        XQ�           .?AVGeModalDialog@@     XQ�           .?AViCustomGui@@        XQ�           .?AVNeighbor@@  XQ�           .?AVC4DThread@@ XQ�           .?AVtype_info@@ u�              2��-�+  �] �f�������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            0  C  �j `  �  �j �  �  pj �  �  xj    N  hj p  ,  �k @  �  �k �  �  �k 0  \   n   <  hk P  |  �k �  �  �j �  C  �j `  �  �j �  �  n �  �  pk �  �  �k �    �j    S  k `  �  k �  �  n    6  xk P  �  �k �    `l    �  �m �  /  �m @  a  �k p  �  �k �  �  `k �  �  �k    $  Xk 0  f   k �  �  Pk �  
  (k    �  �m    s  �j �  B   �m p   �$  �l �%  �)  �m +  �+  dm @,  �,  �m  -  j-  �k �-  �-  8k �-  .  �k 0.  c.  Hk p.  �.  @k �.  m/  �m �/  `0  n p0  �0   n �0  1  (n  1  ?1  0n P1  �1  8n �1  �1  @n 2  >2  Hn P2  j2  Pn p2  �2  Xn P3  h3  �n p3  �3  �n �3  �4  �n �4  A5  o P5  �5  o �5  �5  o  6  �6   o �6  �6  (o �6  18  0o @8  T:  �o `:  <=  Pp P=  A  (q A  _A  0r pA  �A  8r �A  YB  @r `B  D  Hr 0D  BF  �r PF  gF  8s pF  �F  @s �F  �F  `n �F  G  �n G  >G  hn @G  vG  xn �G  �G  pn �G  H  Ps H  �H  Xs �H  �H  Hs �H  (I  �n pI  �I  �s �I  J  �s J  4J  �s @J  �J  �s �J  �J  t  K  *K  t 0K  TK   t `K  zK  (t �K  �K  0t �K  �K  8t  L  $L  @t 0L  JL  Ht PL  ~L  Pt �L  �L  Xt �L  �L  `t  M  M  �t  M  DM  �t PM  �M  �t �M  �M  �t �M  QN  �t `N  �N  u �N  1O  Hu @O  {O  �u �O  �O  �u �O  P  �u  P  AP  �u PP  �P  �u �P  �P  v Q  �Q   v �Q  R  hv 0R  �R  �v �R  �R  �v �R  S   w S  ;S  w PS  {S  w �S  �S  w �S  �S   w T  HT  (w PT  ~T  0w �T  �T  8w �T  �T  @w  U  3U  Hw @U  �U  Pw �U  V  �w V  ;V  �w PV  �V  �w �V  W  �w  W  zW  �w �W  �W   x �W  �W  x �W  X  x 0X  eX  x pX  �X   x �X  �X  (x  Y  !Y  0x 0Y  QY  8x `Y  �Y  @x �Y  �Y  Hx �Y  �Y  Px  Z  .Z  Xx @Z  nZ  `x �Z  �Z  hx �Z  �Z  px  [  .[  xx @[  n[  �x �[  �[  �x �[  �[  �x  \  .\  �x @\  �\  �x �\  ]  �x  ]  ?^  �x P^  �^  (y �^  C_  0y P_  �_  8y �_  }`  @y �`  �`  Hy �`  �`  Py �`  a  Xy 0a  ^a  `y pa  �a  hy �a  �a  py �a   b  xy 0b  `b  �y pb  �b  �y �b  �b  �y �b  Kc  �y `c  �c  �y �c  od  �y �d  �d  �y  e  pe  �y �e  f  �y  f  �f  �y �f  �f   z �f  g  z  g  �g  z �g  h  z h  'h   z 0h  `h  (z ph  �h  0z �h  �h  8z �h  i  @z i  1i  Hz @i  ai  Pz pi  �i  Xz �i  �i  `z �i  j  hz j  �j  pz �j  �j  �z �j  �j  �z  k  !k  �z 0k  Qk  �z `k  �k  �z �k  ul   { �l  �l  h{ �l  �l  p{ �l  m  x{  m  Xm  �{ `m  �m  �{ �m  �m  �{ �m  
n  �{ n  :n  �{ @n  kn  �{ �n  �n  �{ �n  �n  �{ �n  o  �{  o  No  �{ `o  �o  �{ �o  �o  �{ �o  p  �{  p  Mp  �{ `p  �p  �{ �p  �p  �{ �p  �p   | q  ;q  | Pq  {q  | �q  �q  | �q  �q   | r  >r  (| Pr  ~r  0| �r  �r  8| �r  s  @|  s  Ns  H| `s  �s  P| �s  �s  X| �s  t  `| 0t  zt  h| �t  �t  p| �t  �t  x|  u  .u  �| @u  nu  �| �u  �u  �| �u  �u  �|  v  .v  �| @v  nv  �| �v  �v  �| �v  �v  �|  w  .w  �| @w  nw  �| �w  �w  �| �w  �w  �|  x  .x  �| @x  nx  �| �x  �x  �| �x  �x  �|  y  .y   } @y  ny  } �y  �y  } �y  �y  }  z  .z   } @z  xz  (} �z  �z  0} �z  {  8}  {  W{  @} `{  �{  H} �{  �{  P} �{  |  X}  |  N|  `} `|  �|  h} �|  �|  p} �|  }  x} }  H}  �} P}  t}  �} �}  �}  �} �}  �}  �} �}  ~  �} ~  *~  �} 0~  `~  �} p~  �~  �} �~  �~  �} �~  <  �} P  �  �} �  �  �} �  �  �} �  9�  �} @�  u�  �} ��  ��  �} ��  �   ~  �  !�  ~ 0�  �  ~ �  1�  x~ @�  k�  �~ ��  ̂  �~ ��  "�  �~ 0�  T�  �~ `�  ��  �~ ��  �  �~  �  ��  �~ ��  Մ  8 ��  ߅  @ ��  o�  � ��  ��  � ��  ��   �  �  $�  � 0�  ��  � ��  �  X�  �  .�  `� 0�  `�  ht `�  ��  xt ��  ܈  pt ��  �  �t p�  ��  x� ��  �  ��  �  8�  �� @�  n�  �� ��  ��  �� ��  �  �� �  R�  �� `�  ��  �� ��  ߋ  �� ��  5�  �� @�  q�  Ȁ ��  ��  Ѐ ��  ߌ  ؀ ��  )�  �� 0�  W�  � `�  ȍ  �� Ѝ  �  �� ��  .�   � @�  ��  � ��  &�  � 0�  ��  � ��  ��   � ��  �  (�  �  '�  0� 0�  a�  8� p�  ��  @� ��  �  H� �  !�  P� 0�  a�  X� p�  ��  `� ��  ��  h� �  7�  p� @�  g�  x� p�  ��  �� ��  ג  �� ��  �  ��  �  G�  �� P�  w�  �� ��  ��  �� ��  �  ��  �  e�  �� p�  ��  �� ��  ��  ȁ �  K�  Ё `�  ��  ؁ ��  Ε  �� ��  ��  �  �  +�  �� @�  n�  �� ��  ��   � ��  ٖ  � ��  �  � 0�  J�  � P�  ��   � ��  �  (� �  V�  0� `�  ��  8� ��  �  @�  �  Q�  H� `�  ��  P� ��  ֙  p� ��  /�  X� @�  �  `�  �  (�  8� 0�  K�  @� Р  �  H� �  *�  �� 0�  c�  �� p�  ��  �� ��  ޡ  �� �  8�  �� @�  ��  �� ��  ΢  ȃ �  �  Ѓ  �  X�  ؃ `�  ��  �� ��  %�  � 0�  T�  0� `�  ��  8� ��  ��  @� Ф  ��  H� �  *�  P� 0�  J�  X� P�  j�  `� p�  ��  h� ��  ��  p� ��  �  x� �  B�  �� P�  ��  �� ��  Ѧ  �� �  (�  �� 0�  ^�  �� p�  ��  �� ��  �  �� �  \�  � p�  ��  �� ��  �  �� �  W�   � `�  ��  � ��  ��  �  �  ��  � ��  �   �  �  ��  (� ��  ƫ  0� Ы  ��  8� �  4�  @� @�  d�  H� p�  ��  P� ��  ̬  X� �  �  `�  �  D�  h� P�  ��  p� ��  �  x� 0�  F�  �� P�  ��  ȅ ��  �  Ѕ �   �  ؅ 0�  
�  �� �  �  �  �  X�  �� `�  ��  �� ��  ��   � ��  �  �  �  �  �  �  S�  � `�  ��   � ��  Ӳ  X� `�  ѳ  �� �  F�  �� P�  ��  І ��  ݶ  ؆ �  �  ��  �  �  � ��  	�  �� �  ;�  �� P�  q�   � ��  ��  � ��  ֹ  � �  �  �  �  t�   � ��  Ժ  (� �  .�  0� @�  ��  8� ��  7�  @� @�  ��  H� ��  �  P�  �  �  X�  �  `�  �� p�  ɾ  �� о  ��  �� ��  "�  ȇ 0�  ��  Ї ��  ��  ؇  �  U�  �� `�  ��  @� ��  ��  X� ��  @�  p� @�  ��  X�  �  ;�  x� @�  c�  `� ��  ��  � ��  ;�   � @�  ��  � ��  ��  �  �  E�   � P�  ��  �� ��  )�  (� 0�  |�  �� ��  ��  � 0�  T�  h� `�  ��  0� ��  ��  H� ��  @�  �� @�  ��  8� ��  ��  P� ��  �  �� `�  ��  � @�  ��   � ��  ��  (� P�  ��  0� ��  ��  8� ��  '�  p� 0�  U�  x� `�  ��  �� ��  ��  �� ��  ��  �� ��  �  ��  �  M�  �� `�  ��  �� ��  ��  �� ��  �  ��  �  P�  �� `�  ��  ȉ ��  ��  Љ ��  S�  ؉ `�  ��  �� ��  ��  � ��  *�  �� 0�  l�  �� ��  n�   � ��  ��  � ��  �  �  �  f�  � p�  ��   � ��  	�  (� �  ��  0� ��  ��  8� �  u�  @� ��  ��  H�  �  -�  P� @�  o�  X� ��  ��  `� ��  ��  h�  �  (�  p� 0�  d�  x� p�  ��  �� ��  ��  ��  �  (�  �� 0�  |�  �� ��  ��  ��  �  <�  �� P�  ��  �� ��  ��  �� ��  ,�  �� @�  ��  Ȋ ��  #�   � 0�  j�  � p�  ��  � ��   �  � �  h�   � p�  ��  (� ��  C�  0� P�  ��  8� ��  ��  @�  �  (�  H� 0�  X�  P� `�  ��  X� ��  �  `� ��  ��  h� ��  ��  p� ��  �  x� �  ,�  �� @�  D�  �� P�  ��  �� ��  ��  � ��  5�  �� @�  ��  �� ��  ��   � ��  j�  � p�  ��  � ��  ��  �  �  %�   � 0�  ��  (� ��  �  0�  �  ��  8� ��  �  @�  �  ��  �� ��  K�  �� `�  d�  �� p�  �   �  �  Z�  � `�  0�  `� @�  ��  �� ��  c�  �� p�  �  ��  �  ��   � ��  �  �  �  ��  � ��  ��  � ��  -�   � @�  ��  (�  �  ��  4� ��  .�  |� @�  ��  �� ��  �  ��  �  ��  �� ��  9  �� @  �  �� �   ��   � �� � x �� � - � @ � l�   T t� ` � |� �  ��   { �� � # �� 0 � �� � ( ԏ 0 � � �  � 0 � � � x	 $� �	 �	 ,�  
 u
 4� �
 �
 <�   y D� � � L� � � T� � 4 � @ � �� � � ��  \ � p � � �  � 0 � � � > $� P � ,�   j 4� p  <�   � D� � u L� �   T� 0 � \� � � d� � - l� @ � t� � � |� � = �� P � ��   � �� � R �� `  ��  � �� � P �� ` � ��   � đ � 0 ̑ @ � ԑ � � ܑ �   �    �  � �  ~! �� �! " �� " �" � �" -# � @# $ �  $ �$ � �$ #% $� 0% �% ,� �% #& 4� 0& �& <� �& ' D� 0' h' L� p' �' T� �' ( \�  ( `( d� p( �( l� �( �) t� �) g* �� p* �* ��  + �+ �� �+ �+ Ē �+ i, ̒ p, �, Ԓ �, $- ܒ 0- �- � �- >. � P. �. �� �. ^/ �� p/ �/ � 0 �0 � �0 F1 � P1 �1 � �1 U2 $� `2 �2 ,� �2 E3 4� P3 �3 <� �3 B4 D� P4 �4 L� �4 %5 T� 05 �5 \� �5 #6 d� 06 s6 l� �6 t7 t� �7 �7 �� �7 ;8 �� P8 �9 �� �9 R: ē `: 7; ̓ @; h; � p; < �  < �< d� �< 4= �� @= g= Ĕ p= > ̔  > H> Ԕ P> �? ܔ �? 4A � @A �B � C fC �� pC �C �� �C &D � 0D hD � pD �D � �D BE � PE �E $�  F gF \� �F IG d� PG �G �� �G H �� 0H VH �� `H �H ĕ �H I ̕ I �I � �I �I <� �I 2J D� @J �J L� �J zK �� �K �K �� �K �K Ė  L RL ̖ `L �L Ԗ �L M ܖ  M `N $� pN �N �� �N  O �� O 2O �� @O �O ė �O �R ̗ �R �S �� �S �U ܘ  V �W t� �W X ̙ 0X `X ԙ �X Z ܙ 0Z c[ � p[ �[ <� �[ \\ D� p\ R] L� `] j^ Ě p^ �^ � �^ \_ � p_ �_ � �_ _` $� p` �` ,� a Ib 8� Pb �b D� �b �c P� �c  d �  d td �� �e �e � �e �e |� �e f ��  f �f h� �f 2g p� @g |g Ј �g �g ��  h ah Ȉ ph �h d� �h �h l� �h &i \� 0i fi ؈ pi �i t� �i �i �� k �k X� �k l l� l �l � �l �l �� �l �l `�  m 6m �� @m �m  � �m �m h�  n ,n �� @n �n ̛ �n o �� o 1o x� Po �o �� �o �o � �o p H�  p Kp  � Pp {p P� �p �p d� �p �p � �p q � pq �q �� �q �q ě �q r  � Pr �r p� �r �r �� �r s �� s 9s �� @s us x� �s �s �� �s �s ��  t (t � 0t Wt � `t �t �� �t �t �� �t u ȝ u <u Н Pu �u ؝ �u �u �� �u v �  v Gv � Pv v �� �v �v  � �v �v � w Iw � Pw �w � �w �w  � �w x (�  x ox 0� �x �x 8� �x 	y @� y Ay H� Py wy P� �y �y X� �y �z `� �z �z �� �z { ��  { Q{ �� `{ �{ �� �{ �{ �� �{ �{ ��  | �~ Ȟ �~ �~ О   ' ؞ 0 W �� ` � � � � � � � �� � 7�  � @� g� � p� �� � �� � � �� � $�  � O� ,� `� �� 4� �� Ӂ <� �� � D�  � Q� L� `� �� T� �� "� \� 0� N� d� `� �� l� �� ǃ t� Ѓ �� |�  � 1� �� @� o� �� �� �� �� �� �� ��  � =� �� P� � �� � C� �� P� w� �� �� �� ğ �� ׆ ̟ �� � ԟ � 7� ܟ @� y� � �� Ç � Ї � �� 0� �� �� �� )� � 0� !� � 0� W� � `� �� � �� � $�  � '� ,� 0� W� 4� `� �� <� �� э D� �� � L� � A� T� P� w� \� �� �� d� Ў � l� � A� t� P� �� |� �� Ϗ �� �� � ��  � G� �� P� �� �� А � �� � U� �� `� �� �� �� Ǒ �� Б 	� Ġ � -� ̠ @� g� Ԡ p� �� ܠ В �� �  � r� � �� � ��  � '� � 0� i� � p� �� � �� � � � #� $� 0� �� ,� �� ߕ 4� � ?� <� P� �� D� �� ܖ L� � ;� T� P� g� \� p� �� h� �� � p� � t� x� �� � ��  � [� �� p� �� �� �� 6� �� p� �� �� �� C� �� P� �� �� �� �� ��  � d� �� p� �� ȡ Ю !� С 0� � ء  � m� � �� Ͱ � � � � � �� �� б }�  � �� �� � �� � �  � '� � 0� k�  � p� �� �� �� � � � � � � )�  � P� �� �� �� Ե �� � � X� p� �� p�  � �  �  � Q� H� p� �� �� �� � �� � 4� � @� g� �� p� �� �� �� �� h� �� � `� � � �� � -� �� 0� P� �� P� p� �� p� �� x� �� �� p� �� � (� � � @�  � Y� 0� `� �� 8� �� ļ x� м �� Т  � Q� �� `� �� 0� �� � h� � � P� � ;� آ @� q� Ȣ �� �� �� �� &� � 0� s� � �� *� � 0� f� �� p� �� �� �� �� �� �� ?� `� @� � P� � -� @� 0� �� � �� � � 0� �� \� �� �� �� `� �� � �� �� � �� �� �� �� �� ̣  � � �� @� 	� � � �� ��  � �� ԣ �� � �  � �� �� �� � �� � �� �� �� l� �� p� u� �  � p� �� p� �� � �� �� x� �� � t� P� �� (� �� �� 0� �� � �  � D� � P� |� �� �� �� � �� 5� �� @� �� \� �� �� D� �� � l�  � X� d� `� z� �� �� �� P� ��  � 8�  � Y� |� `� �� �� �� �� �� � o� �� �� �� �� �� O� �� `� �� �� �� g� �� p� �� �� �� � ĥ  � p� ̥ �� �� ԥ �� %� ܥ 0� �� � �� �� � �� _� �� p� 9� �� @� �� T� �� �� \�  � ;� d� P� � l�  � �� t� �� W� |� �� �� Ԧ �� � ܦ  � �� � �� �� � �� ,� �� @� �� �� �� �� � �� @� � P� �� � �� � �  � b� $� p� �� ,� �� *  4� 0  s  <� �  �  D� �   L�   u T� � � \� �  d�   c l� p � t� � ' |� 0 � �� � � �� � 1 �� @   �� 0 � �� � � ��   R � ` � � �  �  v � � � $� � F ,� P � 4� � 	 <� 	 �	 D� �	 �	 �� 0
 �
 �� �
 � �� � � ��   @ � P r � � � �   V � ` � $� � � ,�   _ 4� ` � <� � � D� � � L� �  T�   N l� ` � t� � � |� � � ��   - �� @ k �� � � �� �   ��  @ �� P  �� � � �� �  ĩ   N ̩ P � ԩ � � ܩ � � \�   / d� 0 \ � ` � � � � �� � � ��  ' � 0 c � p � � �  � 0 F $� P � ,� � � 4� �  <�   A D� P { L� � � T� � % \� 0 o d� � � l� �  t�  O |� ` � �� �  �� 0 J �� P j �� p � �� � � ��  w �� � � �� � � � � � �    �   X � ` � $� � � ,� � � 4�   Q <� ` � D� � 
 L�  H �� P t �� � � ��    n  �� �  �  D� �  �  L� ! :! T� @! j! \� p! �! d� �! �! l� �! �! t�  " $" |� 0" J" �� P" r" �� �" �" �� �" �" �� �" �" �� �" # ��  # T# �� `# �# �� �# �# Ĭ �# $ ̬  $ L$ Ԭ `$ �$ ܬ �$ % $�  % b% ,� p% �% 4� �% �% <� �% 
& D� & z& L� �& �& �� �& �& �� �& ' ��  ' L' �� `' �' �� �' �' �� �' &( ȭ 0( f( Э p( �( ح �( �( � �( ) �  ) L) � `) z) �� �) �)  � �) * � 0* R* � `* �* � �* �*  � �* 6+ (� @+ �+ p� �+ �+ �� �+ , ��  , _, Ȯ p, �, Ю �,  - خ - D- � P- z- � �- �- � �- �- �� �- .  � . 4. � @. l. � �. �. � �. //  � @/ d/ h� p/ �/ p� �/ �/ x� �/ �/ �� �/ �0 �� �0 �0 �� �0 |1 �� �1 ,2 �� @2 �2 �� �2 �2 ��  3 63 �� @3 �3 ȯ �3 �3 Я �3 4 د 04 J4 � P4 �4 � �4 5 �  5 �5 8�  6 $6 �� 06 �6 �� �6 7 ��  7 �7 Ȱ �7 8 � �8 9 X�  9 : �� : �: �  ; �; �� �; 7< ز @< �< 0� �< �< 8�  = 8= @� @= ~= H� �= �= P� �= �= X� �= (> `� 0> h> h� p> �> p� �> �> x� �> 
? �� ? q? �� �? �? �� �? @ �� @ *@ �� 0@ f@ �� p@ �@ �� �@ �@ �� �@ &A �� 0A TA � `A �A � �A �A � �A �A  �  B 6B (� @B xB 0� �B �B 8� �B �B @�  C $C H� 0C \C P� pC �C X� �C �C `� �C �C h� �C 
D p� D xD x� �D �D �� �D �D �� �D E �� 0E �E �� �E EH �� PH �H �� �H J �� 0J �J ȴ �J FK д PK jK �� �K �K �� �K �K ش  L L � 0L �L � �L �L � �L =M �� PM �M  � �M �M �  N |N � �N P �  P ^P  � pP +Q (� @Q jQ 0� pQ �Q 8� �Q �Q @� �Q �Q H�  R 'R P� 0R MR X� `R �R `� �R �R h� �R �R p� S 7S ȵ @S {S е �S T ص T 7T � @T {T � �T �T � �T �T �� �T U  �  U SU � `U �U � �U &V X� 0V _V `� pV �V h� �V �V p� �V �V x�  W BW �� PW �W �� �W �W �� �W *X �� 0X TX �� `X �X �� �X �X �� �X �X �� �X +Y �� @Y {Y ȶ �Y �Y ж �Y -Z ض @Z qZ � �Z �Z � �Z �Z �  [ ;[ �� P[ �[  � �[ �[ � �[ \ � 0\ k\ � �\ �\  � �\ �\ (� �\ $] 0� 0] g] 8� p] �] @� �] �] H� �] ^ P�  ^ �^ X� �^ o_ �� �_ �_ �  ` �` `� a b ظ  b �b P� �b c ��  c �c  � �c kd h� �d ?e �� Pe �e (� �e �f �� �f 9g � @g $h D� 0h �h �� �h 	i � i fi � pi Tj  � `j �j �� �j �k � �k Il P� Pl m ��  m �m � �m �n h� �n 	o Կ o �o ,� �o Wp �� `p q �� 0q �q T� �q r �� r 7r �� @r gr �� pr �r �� �r �r ��  s /s �� @s gs �� ps �s �� �s �u �� �u �u \�  v 'v d� 0v _v l� pv �v t� �v �v |� �v �v �� w *w �� 0w cw �� pw �w �� �w �w �� �w 'x �� 0x ux �� �x �x �� �x %y �� 0y �y �� �y �y �� �y �y ��  z /z �� @z {z �� �z �z �� �z { �� 0{ k{ � �{ �{ � �{ �{ � �{ �| � �| �| $� �| 
} ,� } 4} 4� @} d} <� p} �} D� �} �} L� �} k~ T� �~ �~ \� �~ 2 d� @ q l� � � t� �  |� Ѐ �� �� �� � \� �� !� d� 0� M� l� `� }� t� �� �� |� �� � �� �� "� �� 0� t� �� �� �� �� �� � �� �� ;� x� �� � �� `� }� �� ��  �� Ѕ �� ��  � /� �� 0� W� �� `� �� �� �� �� �� �� � �� �� � ��  � C� �� P� �� �� �� �� �� �� � �� �� � ��  � D� �� P� y� �� �� �� �� �� � �� �� � �  � D� � P� t� � �� �� � �� � $� �� � ,�  � D� 4� P� t� <� �� �� D� �� Ԋ L� �� � T� � 4� \� @� c� d� p� �� l� �� ԋ t� �� � |� � 6� �� @� s� �� �� �� �� �� Ԍ �� �� � �� � C� �� P� �� �� �� � �� �� 6� �� @� �� �� �� Ύ �� �� � ��  � N� �� `� �� �� �� ̏ � �� � �  � @� � P� �� � �� �� $� �� � ,� � (� 4� 0� T� <� `� �� D� �� � L� � � T�  � S� \� `� �� d� В � l�  � 3� t� p� �� |� �� ē �� Г �� �� � F� �� P� |� �� �� �� �� �� � ��  � 6� �� @� �� �� �� Ε �� �� � ��  � Q� �� `� �� �� �� Ė �� Ж � �� � <� �� P� � �� � �� � �� ɘ � И � � � �� $� �� �� 4� �� ٚ <� �� �� D�  � �� L� �� � \� � /� d� 0� 4� l� �� �� �� �� D� �� P� �� �� �� ן �� �� ؠ �� � $� �� 0� �� �� �� ~� �� Ф �� �� �� ʬ �� Ь �� �� ��  � �� � �� �� �� �  �  � �� � �� 	� � � �� � �� �  �  � �� (� �� �� 0� �� � 8�  � Z� @� `� �� H� �� � P�  � �� X� �� ܷ `� � <� h� P� �� p� �� � x� � 2� �� @� �� �� �� � �� � 2� �� @� �� �� �� ں �� � 2� �� @� �� �� �� � �� � 8� �� @� �� �� �� ּ �� � &� �� 0� �� �� �� � ��  � v� �� �� �  � � L� � `� �� � �� � � 0� ��  � �� �� (�  � �� 0� �� .� 8� @� �� @� �� � H�  � p� P� �� �� X� �� D� `� �� � h� � C� �� P� �� x� �� \� �� `� �� �� � \� �� �� �� �� �� �� p� �� !� �� 0� d� �� p� �� �� �� � �� 0� r� �� �� �� �� �� � �� 0� m� �� �� �� �� �� � ��  � �� �� �� g� �� p� � �  � o� p� �� �� x� �� �� �� �� $� �� 0� �� �� �� �� �� �� �� �� �� �� �� � {� �� �� �� �� �� 	� �� � I� �� P� �� �� �� =� �� P� �� �� �� '� �� 0� }� �� �� �� �� �� �  �  � k� � �� �� � �� %� � 0� v�  � �� 9� (� @� � x� � 8� �� @� �� �� �� �� �� �� � �� 0� �� �� �� � �� � q�  � �� �� X� �� b� 0� �� '� h� 0� �� x� �� w� p� �� �� �� �� 1� �� P� 1� �� @� �� ��  � 3� �� P� �� � �� ��  � �� �� �  � K� ,� P� !� 4� 0� C� $� P� �� � �� �� � � �� <� �� �� �� �� @� d� `� � �� � �� �� �� � ��  � 2� �� @� ~� �� �� �� �� �� �� �� �� �� 8l �� �� @l �� ˶ Hl � � �l  � 8�  k 8� ^� k p� �� Dm �� �� Lm �� �� Tm �� ܷ \m  � � �m � 0� �m @� X� �n X� ��  o �� �� �o �� �� �o �� ݸ �o ݸ �� 0p �� � 8p � 6� @p 6� Q� Hp Q� i�  q i� �� q �� �� q �� ¹ q ¹ ݹ  q ݹ ��  r �� � r � 6� r 6� Q� r Q� l�  r l� �� (r �� �� �r �� ˺ �r ˺ �� �r �� �  s � 8� (s 8� a� 0s p� �� �s �� �� �s �� Ȼ  t Ȼ � t  � � �t � 0� u 0� H� @u H� `� xu `� x� �u x� �� v �� �� v �� μ Xv μ �� `v �� � �v � 8� �v 8� P� �v P� y� �v y� �� �w �� �� �w �� Ͻ �w Ͻ �� �w �� � �x � %�  y %� =� �y =� U� �z U� ~� �z ~� �� { �� �� { �� ׾ X{ ׾ �� `{ �� � p~ � -� �~ -� V� �~ V� n� ( n� �� 0 �� �� � �� � � � � � � '� � '� P� � P� h� H� h� �� P� �� �� � �� �� � �� �� � �� ��  � �� � (� � /� 0� 0� H�  � H� n� (� n� �� �� �� �� �� �� �� �� �� �� P� �� �� �� �� (� Ȇ (� @� �� @� X� �� `� x� h� x� �� �� �� �� Ћ �� �� ؋ �� �� �� �� � �� � � �� � 1� � 1� I� P� I� a� X� a� y� �� y� �� �� �� �� �� �� �� t� �� �� � �� �� � �� 	� \� 	� !� d� !� 9� ̏ 9� Q� � Q� i� ̐ i� �� Ԑ �� �� ܐ �� �� � �� �� �� �� �� �� �� �� �� �� � T� � )� \� )� A� �� A� Y� �� Y� q� T� q� �� �� �� �� �� �� �� �� �� �� 4� �� �� |� �� � �� � '� � '� M� � M� e� �� e� }� �� }� �� �� �� �� �� �� �� t� �� �� |� �� � �� � *� �� *� E� �� E� `� �� `� x� Ԙ x� �� T� �� �� \� �� �� d� �� �� l� �� �� �� �� � ę � )� 4� )� A� �� A� Y� �� Y� t� �� t� �� � �� �� ؜ �� �� �� �� �� �� �� � �� � (� @� 0� H� X� H� n� `� p� �� � �� �� � �� �� �� �� �� T� �� � �� � +� ؤ 0� V� D� V� n� L� n� �� Ħ �� �� ̦ �� �� � �� �� � �� � �� � +� �� 0� K� �� P� h� � h� �� �� �� �� �� �� �� �� �� �� � �� �� �� �� � 4� � :� <� :� R� � R� x� � x� �� �� �� �� �� �� �� `� �� �� h� �� � �� � 2� �� 2� J� X� J� s� `� s� �� (� �� �� 0� �� �� �� �� �� �� �� 
� �� 
� "�  � "� K� � K� c� H� c� �� P� �� �� �� �� �� � �� �� �� �� ��  � �� #� h� #� ;� p� ;� S� x� S� k� Ȳ k� �� в �� ��  � �� �� (� �� �� �� �� ��  �  � � H� � >� P� >� V� �� V� |� �� |� �� �� �� ��  � �� �� P� �� �� X� �� �� �� �� � ȸ � 5� и 5� M� 8� M� e� @� e� �� H� �� �� �� �� �� �� �� �� � �� �� �� �� � X� � � `� � 6� �� 6� N� �� N� f� � f� ~�  � ~� �� p� �� �� x� �� �� ܻ �� �� � �� �� 4� �� � <� � &� �� &� >� �� >� V� �� V� n�  � n� �� |� �� �� �� �� �� Խ �� �� ܽ �� �� @� �� �� H� �� � �� � .� �� .� F�  � F� ^� � ^� v� X� v� �� `� �� �� Ŀ �� �� ̿ �� �� � �� �� $� �� � �� � � �� � 6� �� 6� N� �� N� f� D� f� ~� L� ~� �� �� �� �� �� �� �� L� �� �� T� �� �� �� �� � �� � )� L� )� A� T� P� h� X� h� �� `� �� �� h� �� �� �� �� �� �� �� � �� � *� �� *� E� �� E� `� �� `� {� �� {� �� �� �� �� �� �� �� � �� �� P� �� � h� � 1� p� @� p� �� p� �� �� �� �� �� �� �� \� �� � �� � M� �� �� �� �j �� �� �k  � !� �s 0� L� h� P� l� P� p� �� �� �� �� �� �� �� �� �� ��  � �� � �� � ,� �� 0� D� |� P� �� t� �� �� � �� �� `� P e �s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �`         f `c @`         �h �b                         Rh     <h     "h     h     �g     �g     �g     hh                                                                                                     �e     �e     �e     �e     �e     �e     �e     �e     �e     �e     f     (f     6f     Df     Pf     df     �e     ~f     �f     �f     �f     �f     �f     �f     �f     �f     g     (g     Fg     dg     xg     �g     �e     �e     |e     re     he     `e     Ve     pf     @e                                                                                                                                                             Rh     <h     "h     h     �g     �g     �g     hh                                                                                                     �e     �e     �e     �e     �e     �e     �e     �e     �e     �e     f     (f     6f     Df     Pf     df     �e     ~f     �f     �f     �f     �f     �f     �f     �f     �f     g     (g     Fg     dg     xg     �g     �e     �e     |e     re     he     `e     Ve     pf     @e                                                                                                                                                             �__CxxFrameHandler3  =memset  �free  .malloc  ;memmove �floor 9memcpy  pstrlen  �asin  �cos `sqrt  �fabs  �fmod  1_purecall 	_vsnprintf  ostrftime  z_localtime64  �_time64 jstrcpy  MSVCR110D.dll �__CppXcptFilter _amsg_exit  �_malloc_dbg �_free_dbg __CrtSetCheckCount _initterm _initterm_e �__C_specific_handler  |_lock �_unlock N_CrtDbgReportW  2_calloc_dbg �__dllonexit %_onexit �__crt_debugger_hook �__crtUnhandledException �__crtTerminateProcess �__crtCaptureCurrentContext  �__crtCapturePreviousContext :?terminate@@YAXXZ "?_type_info_dtor_internal_method@type_info@@QEAAXXZ �__clean_type_info_names_internal  �IsDebuggerPresent @EncodePointer DecodePointer �IsProcessorFeaturePresent ?QueryPerformanceCounter *GetCurrentProcessId .GetCurrentThreadId  �GetSystemTimeAsFileTime KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                     �   � �0�8�@�H�P�X�`�h�p�x�������Ф������ ���� �(�0�8�@�H�P�X�`�h���������������ȪЪت����� ���� �(�0�8�@�H�P�X�`�h�p�x�������������� ���� �(�0�8�@�H�P�X�`�h�p�x�������������������ȬЬج�謰���   0 |   0�8�@�H�P�X�`�h�p�x�������������������ȮЮخ����� ���� �(�0�8�@�H�P�X�`�h�p�x�������������������ȯЯد����� @ $    ���� �(�������� �(�0�8� P    P�X�� ���   �      �(�P�x���Ƞ��8�`�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                