MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       "�r8f�kf�kf�ko܏ke�kf�k,�k��kg�k	҂kx�k	Ҷk
�k	ҷk^�k	҇kg�k	ҁkg�kRichf�k                PE  L �pQ        � !
  �  �      ��     �                       �         @                   @ H   t (                            ` �                                  � @            �                           .text   O�     �                   `.rdata  �Z   �  \   �             @  @.data   �1                      @  �.reloc  �"   `  $   "             @  B                                                                                                                                                                                                                                                                                                                                                                                                �  �   �����̋D$Ht�   ù`3�  ������������������������̡p3V��H�QV�ҡp3�T$�H�D$�IRj�PV�у���^� �����������̡p3�P�BQ��Y�V�t$W3���t.S�\$U�l$SU����  �p3���   �B(��G�Ћ���u�][��_^��V�t$W3���t?S�\$U�l$�D$P���~  ;�uG��u�p3���   �B(���Ћ���u�][��_^Ë�_^Ã�$�p3�H�A�T$VR�Ћp3�Q�Jj j��D$h��P�у��T$R�L$��+  �p3�H�A�T$R�Ћp3�Q�J�D$P�ыp3�B�Pj j��L$(h��Q�ҋD$��j P�L$ Qh@ j j �  ��PhD� �A@  �p3���B�P�L$4Q�҃� �L$�,  ��^��$���������������P�X�����D$����D$�X�D$�X� ������̡p3V��H�QV�҃���^��������̡p3V��H�QV�ҡp3�H�T$�AVR�Ѓ���^� ��̡p3�H�T$�I(��VWR�D$P�ыp3�t$$���B�HV�ыp3�B�HVW�ыp3�B�P�L$Q�҃�_��^���̡p3�P���   ��p3�P�D$���   ��P�D$$P�D$P�ҋL$���P�Q�P�Q�P�Q�P�@�Q�A����� �p3�P�R4����̡p3�P�RH����̡p3�P�R8����̡p3�P@�B,Q�Ѓ���������������̡p3�P�BQ�Ѓ���������������̡p3�P�BQ�Ѓ���������������̃�HV�t$TW������? HP����D � /�������   S�$�� �|$Xjj?��� P�x��������  �p3�H@�Q,W�ҋ��p3�H�A(�T$ VR�Ћp3�Q�J���D$P�ыp3�B�P�L$QV�ҡp3�H�A�T$4R�Ћp3�Q�R8���D$PS���ҡp3�H�A�T$R�Ѓ�[_^��H� �|$Xjj?��3��� P��������G����p3���   �|$X�B4����jj?P���������  �����p3���   �|$X�B4jj?��3���P�h�������  ������L$���  �L$8jQ�6�  ��P�L$ ���  �L$8���  �p3�B�P�L$Q�҃��D$Pj��  ��Pj j�L$,���  �p3�Q�J���D$P�у�����   �O�w��u	�O  ���P  ���u"j�  P貵  ���L$�F�  [_^��H� j j��T$$R��P  ��t"j裵  V��N  ���L$��  [_^��H� �N  j j��j@j@���bP  �jjh   W�R  V�N  ���>�L$���  [_^��H� � �G�5���P�N  ��[_^��H� ��  �  � � � 5 l �p3�H@�Q,�� SUVW�|$4W�҃��ϋ��� ��3ۅ�t*�I j?���  ��uC�p3���   �B(���Ћ���uًp3�Q�J(�D$ SP�ыp3���B�P�L$Q�ҡp3�H�A�T$RV�Ћp3�Q�J�D$4P�ыp3�B�P8���L$Qh�  ���ҡp3�H�A�T$R�Ћp3���   �B4�����Ћ�3���t(j?����  ��uG�p3���   �B(���Ћ���u؋p3�Q�J(�D$ WP�ыp3���B�P�L$Q�ҡp3�H�A�T$RV�Ћp3�Q�J�D$4P�ыp3�B�P8���L$Qh�  ���ҡp3�H�A�T$R�Ѓ�_^][�� � ���������̃�X�IS�\$dUVW�;�73�|$4;�t@;�tV�JM  ��#M  ��p3�H�QV�l$ �l$$�҉D$�p3�H�QV�҃��K;�u�L  Uj��j@j@����M  WhD� � N ����t�V��L  �G�O�W�D$�G�L$ �T$�D$;��x  �p3�Q@�D$l�J,P�ыp3���؋B���   Uh�  ���ҋ���
  ��p3�T$8�L$P�T$@�\$H�P���   �D$8Ph�  Q����� �@�@�P�������� ���ʉD$0��� �ɉD$,��� �ΉD$(��O  �؋D$�L$l�������ŉD$�p3���   �B4�Ћ����   ��I j?���w  ��t�p3���   �B(���Ћ��u��}   3�9l$~u�|$|g�L$�T$ �D$�|��D$$��p3�Q�D$(�L$,P�D$4Q��  PWUV�у���t�p3�B��  h�   WUSV�у�O�L$$u��|$4E;l$|��L$l��  �����   �d$ j?���  ��t�p3���   �P(���ҋ��u��|   3�9l$~t�|$|f�D$�L$�T$�|��T$l��p3�H�T$(�D$,R�T$4P��  RUWV�Ѓ���t�p3�Q��  h�   UWSV�Ѓ�O�L$lu��|$4E;l$|��L$�T$ �D$�O�L$�W�T$p�7�G�O_^]�B   [��X� _^�k][��X� �������̃�SV�t$$WV����  �؅�u	_^[��� �p3�H@�Q,V�ҋ�p3�P�B4��jh�  �����h��p3�\$��D$�\$P�X�h�  �\$$�Q�RH���҃ �Gt	P��H  ��_^��[��� ����̋D$VP���S  �~ �F^tP�H  Y� ��������������̋D$S�\$VWP��L$SQ���E  ����u_^3�[� �T$R�����  ��t�N��t��I  ��$H  �F�|$ t�FP����  ��t���_^[� ��̋D$SVW�|$WP����  �؅�u_^3�[� 3�9N��Q�����  ��t�v��tjj h�� V����  ��t�_^��[� ������S�\$U�l$VW�|$SUW���  �D$��u_^][� ��t4��t���F u0SW��������D$_^][� W�������D$_^][� SW���%����D$_^][� ���������̋D$�T$SV�t$WP�D$���L$ QRPV����  �؅�u_^[� ���> t	V�G  ���O�G  _�^��[� ������������V���  �D$t	V�$  ����^� ��Vhp�j>h�3j�l%  ������t���L  �����^�3�^���������������U��Q�} t�E�E���`3�� �E��M�Q�UR�EP� 6 ����]����������U��Q�M��E��     �M��A    �U��B    �E��@    �E���]������������U��Q�M��M��   ��]��������������U����M�E�x t�o�M�9 t �U�P�p3�Q<�B�Ѓ��M��    �U�z t>�E�x t+�M�Q�U��E��E��}� tj�M��
  �E���E�    �M��A    ��]����������U���$�M܍E�P�>�  ��P�M��   �E��M��W�  �E���]�U����M��E��x uMh��j;h�3j�#  ���E��}� t�MQ�M����  �E���E�    �U��E�B�M��y u3��G�U��z t�E�3Ƀ8 �����/�UR�p3�H<��҃��M���U��B   �E�3Ƀ8 ������]� ����U��Q�M��E��@   �p3�Q<�B�ЋM���U�3��: ����]��������������U��Q�M��E��x t�   �*�M��y u3���U��BP�M��R�p3�H<�Q�҃���]������������U��Q�M��E��8 u�p3�Q���EP�M��R�p3�H<�Q�҃���]� ����U��`3����]��U��EP�`3����]��������������U���(�EP�`3�|���P�M�����j h���M�����j �M�Q�U�R�M��  ������E�M������E��t�M�@����M������E�9j�M�Q�M��  j�j��UR�E�P�M��  �M�Q�M�%����M��M����E��]�������U���<�EP�`3�����P�M������j h���M������j �M�Q�U�R�M���  ������E�M�������E��t�M�����M�������E�   j�M�Q�M���  j�j��UR�E�P�M���  j h���M��_���j �M�Q�U�R�M��}  ������E׍M��{����Eׅ�t�M�����M��c����E�9j�M�Q�M��p  j�j��UR�E�P�M��  �M�Q�M� ����M��(����E��]��U���P�EP�`3����P�M������j h���M�����j �M�Q�U�R�M���  ������E�M�������E��t�M�p����M������E�   j�M�Q�M���  j�j��UR�E�P�M���  j h���M��?���j �M�Q�U�R�M��]  ������E׍M��[����Eׅ�t�M������M��C����E�   j�M�Q�M��M  j�j��UR�E�P�M��i  j h���M������j �M�Q�U�R�M���  ������EÍM�������EÅ�t�M�����M�������E�9j�M�Q�M���  j�j��UR�E�P�M���  �M�Q�M�k����M������E��]�������������U���d�EP�`3����P�M��3���j h���M�����j �M�Q�U�R�M��2  ������E�M��0����E��t�M������M������E�  j�M�Q�M��"  j�j��UR�E�P�M��>  j h���M�����j �M�Q�U�R�M��  ������E׍M������Eׅ�t�M�[����M������E�   j�M�Q�M��  j�j��UR�E�P�M���  j h���M��*���j �M�Q�U�R�M��H  ������EÍM��F����EÅ�t�M������M��.����E�   j�M�Q�M��8  j�j��UR�E�P�M��T  j h���M�����j �M�Q�U�R�M���  ������E��M�������E���t�M�q����M������E�9j�M�Q�M���  j�j��UR�E�P�M���  �M�Q�M�V����M��~����E��]��������U��EP�p3�Q<�B�Ѓ�]�������U���X�E�    j h���M������P�������E��M�� ����}� u3���   �E�    �E�P�M��@ �M�Q�U�R�M�� A ����   �}���   �M��  �E�}� t7�EP�M��q����M�Pj�M�Q�M��  �M����#  ��t	�E�   ��E�    �U��UӋE���t�e���M��u����M���t�e���M��a����UӅ�t�E��E���L����E��]������U���T�E�    �} u0j h���M������P�������E�M��
����} u3���   �E�    �EP�M��? �M�Q�U�R�M���? ����   �}���   �M��  �E�}� t7�EP�M��[����M�Pj�M�Q�M��  �M����  ��t	�E�   ��E�    �U��U׋E���t�e���M��_����M���t�e���M��K����Uׅ�t�E��E��2�+�}�u%�}� t�MQ�M��q  ���  ��t�U��U�������E��]���U����} u3��   �EP�M��> �E�    �E�    �M�Q�U�R�M���> ��tT�}�t�}�u"�EP�M��w  P��������t�   �*�$�}�u�MQ�M���  ����   ��t�   ��3���]������U��p3�H<�Q��]���������������U��Q�M��M����  �E��t�M�Q�  ���E���]� ����U��Q�M��EP�MQ�UR�p3�P�M��B@�Ћ�]� �������U��Q�M��EP�MQ�p3�B�M��PH�ҋ�]� ����������U��Q�M��EP�MQ�UR�EP�p3�Q�M��BL�Ћ�]� ��U��Q�M��EP�M��   �������]� U��Q�M��EP�p3�Q�M��Bx�Ћ�]� ��������������U��Q�M��E�P�p3���   �BT�Ѓ���]��������������U����M�EP�MQ�U�R�p3�P�M싂�   ��P�M�����M�������E��]� ��������������U��Q�M��E�P�p3���   �BH�Ѓ���]��������������U��E�p3�p3�]������������U��Q�M��E��@    �M��    �U��B    �E��@   �E���]������������U��Q�M��} u�4�} t�EP�M�
  � �} t�MQ�M�
  ��U�R�M�
  ��]� �������U��Q�M��EP�p3�Q@�M��Bd�Ћ�]� ��������������U��Q�M��EP�p3�Q@�M��Bh�Ћ�]� ��������������U��Q�M��EP�MQ�p3�B@�M��Pl�ҋ�]� ����������U��Q�M��EP�MQ�p3�B@�M����   �ҋ�]� �������U��Q�M��EP�p3���   �M����   �Ћ�]� ��������U��Q�M��EP�MQ�p3���   �M����   �ҋ�]� ����U��Q�M��p3�P@�M��Bt�Ћ�]������U��Q�M��p3�P@�M��Bx�Ћ�]������U��Q�M��EP�p3�Q@�M��B|�Ћ�]� ��������������U��Q�M��p3�P@�M����   �Ћ�]���U��Q�M��p3���   �M��Bt�Ћ�]���U��Q�M��EP�p3�Q@�M����   �Ћ�]� �����������U��Q�M��p3�P@�M����   �Ћ�]���U��Q�M��EP�p3�Q@�M����   �Ћ�]� �����������U��Q�M��EP�MQ�UR�EP�p3�Q@�M����   �Ћ�]� ���������������U��Q�M��EP�MQ�UR�p3�P@�M����   �Ћ�]� ����U��Q�M��EP�MQ�UR�p3�P@�M����   �Ћ�]� ����U��Q�M��EP�MQ�p3�B@�M����   �ҋ�]� �������U��Q�M��EP�MQ�p3�B@�M����   �ҋ�]� �������U����M��E�P�p3�Q@�B�Ѓ��E��M�#Mt�U��#U��U��	�E�E�E��M�Q�U�R�p3�H@�Q�҃���]� ���U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��Q�M��EP�M�Q�p3�B@�HL�у���]� ����������U��Q�M��E�P�p3�Q@�BH�Ѓ���]�U��Q�M��EP�MQ�UR�E�P�p3�Q@�B�Ѓ���]� ��U��Q�M��EP�M�Q�p3�B@�H�у���]� ����������U��Q�M��EP�MQ�U�R�p3�H@�Q�҃���]� �������U��Q�M��EP�M�Q�p3�B@�H �у���]� ����������U��Q�M��EP�MQ�p3���   �M��P�ҋ�]� �������U��Q�M��EP�MQ�UR�p3���   �M��B�Ћ�]� ����U��Q�M��EP�MQ�UR�p3���   �M��B �Ћ�]� ����U��Q�M��EP�MQ�UR�EP�p3���   �M����   �Ћ�]� ������������U��Q�M��EP�MQ�UR�p3���   �M���D  �Ћ�]� �U��Q�M��E P���E�$�MQ�UR�EP�MQ�p3���   �M����   �ҋ�]� ���������������U��Q�M��EP�MQ�UR�EP�MQ�p3���   �M����   �ҋ�]� ��������U��Q�M��p3���   �M��B$�Ћ�]���U��p3�H@�Q0��]���������������U��j�EPj �p3�Q@�B4�Ѓ�]���U��j�EPh   @�p3�Q@�B4�Ѓ�]����������������U��EP�MQj �p3�B@�H4�у�]�U��p3�H|���]����������������U��E�8 t�M�R�p3�H|�Q�҃��E�     ]�����U��p3�H|�Q ��]���������������U��E�8 t�M�R�p3�H|�Q(�҃��E�     ]�����U��p3�H@�Q0��]���������������U��E�8 t�M�R�p3�H@�Q�҃��E�     ]�����U��EP�p3�Q@���   �Ѓ�]����U��E�8 t�M�R�p3�H@�Q�҃��E�     ]�����U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��Q�M��EP�M�Q�p3�BH��d  �у���]� �������U��EP�MQ�UR�EP�p3�Q �BH�Ѓ�]�����������U��Q�}qF t�1�E�E��}� u�#�MQ�M��w  �U�R�EP�M�������  ��]�������������U��Q�M��p3�P@�M��BT�Ћ�]������U��Q�M��EP�p3�Q@�M��BX�Ћ�]� ��������������U��Q�M��EP�MQ�p3�B@�M��P\�ҋ�]� ����������U��Q�M��p3�P@�M��B`�Ћ�]������U��EP�MQ�p3�B��T  �у�]����������������U��h��hE  �M�������4 Ph��hE  �M�q�������3 P�p3�H��T  �҃�]�����U��Q�M��EP�p3���   �M��B@�Ћ�]� �����������U��Q�M��EP�p3���   �M��BD�Ћ�]� �����������U��Q�M��EP�MQ�p3�B�M��Pp�ҋ�]� ����������U��Q�M��E�� ���E���]����������U��Q�M��E�� ����]�������������U����M��E��E��}� t,�M��M�U�U��}� tj�E���M���ЉE���E�    �E�    ��]�����U��Q�M��p3�P�M���  �Ћ�]���U��Q�M��p3�P�M���(  �Ћ�]���U��� �M��E�P�p3�Q�M���   ��P�M�6�  �M��~�  �E��]� �����U��Q�M��p3�P�M���$  �Ћ�]���U��EP�MQ�p3�B��  �у�]����������������U��EP�p3�Q���  �Ѓ�]����U��p3�H��  ��]������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�p3�B��x  �у�]����������������U��EP�p3�Q��|  �Ѓ�]����U��p3�H��d  ��]������������U��EP�MQ�p3�B��p  �у�]����������������U��EP�MQ�p3�B��t  �у�]����������������U��Q�M��M��q����E��t�M�Q�p  ���E���]� ����U��Q�M��   ��]� ��������������U��Q�M���]� ���U��Q�M��   ��]� ��������������U��Q�M��   ��]� ��������������U��Q�M��   ��]� ��������������U��Q�M��   ��]� ��������������U��Q�M���]� ���U��Q�M�3���]� �U��Q�M�3���]� �U��Q�M�3���]� �U��Q�M�3���]� �U��Q�M�3���]� �U��Q�M�3���]� �U��Q�M��   ��]� ��������������U��Q�M��   ��]� ��������������U��Q�M��   ��]� ��������������U��E�M�H4�U�B�7 �E�@8 ? �M�A<`? �U�B@�? �E�@D�> �M�AHp? �U�BL0? �E�@P�> �M�Al@? �U�BX�? �E�@\ ? �M�A`�? �U�BdP? �E�@T�? �M�Ah�? �U�Bp�> �E�@t? �M�U�Q �E�M��U�E�B0�M�U�Q(�E�@,    ]������������U���   j h�   ��`���P�  ��j �MQ�UR�EP�MQ��`���R��������E �E�h�   ��`���Q�UR�EPj��5 ����]���������U���   ��\����l'  ��\������\����: u��   �EP�M����  j h ��M�����P�M���  j j��M�Q�U�R�E�P�;�  ��P��|���Q���  ��P��`���R��  ��P��\������(  ������؈E���`����#�  ��|�����  �M���  �M���  �M��P����M����  �M���t��\���R�&  ����\�����]� �����U��Q�M��EP��5  ���M���E���]� ���������������U��Q�M��E�P�`&  ����]����������U��EP�M���   Q�UR�&� ��]�̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U��E�8 t�M�R�p3�H��҃��E�     ]������U��hﾭޡp3�H��@  �҃�]����U��} t�EP�p3�Q��@  �Ѓ�]��������������U��EP�MQ�p3�B���  �у�]����������������U��EP�MQ�p3�B��  �у�]����������������U��p3�H��   ��]������������U��} t�E�x��u�   �3�]����U��Q�=p3 t3�}s	�E�   ��E�E�j j �M�Q�p3�B���   �у��j�UR�   ����]���������������U��Q�}s�E   �E��P��� ���E��}� u3��:�} t�M��Qj �U�R�[� ���E�� �����M����M��t3   �E���]������U��Q�=p3 t3�}s	�E�   ��E�E�j j �M�Q�p3�B���   �у��j�UR�E�������]���������������U��Q�=p3 t3�}s	�E�   ��E�E�j j �M�Q�p3�B���   �у��j�UR���������]���������������U��Q�=p3 t3�}s	�E�   ��E�E�j j �M�Q�p3�B���   �у��j�UR��������]���������������U��Q�} t=�E�E��=t3 t�M�y��u�U��R�� ����E�P�p3�Q��Ѓ���]������U��Q�} t=�E�E��=t3 t�M�y��u�U��R蠹 ����E�P�p3�Q��Ѓ���]������U��EP�p3�Q��Ѓ�]��������U��EP�p3�Q��Ѓ�]��������U��Q�=p3 t7�}s	�E�   ��E�E��MQ�UR�E�P�p3�Q���   �Ѓ��j�MQ�A�������]�����������U����=p3 tv�} t9�}s	�E�   ��E�E��MQ�UR�E�P�p3�Q���   �Ѓ��I�7�}s	�E�   ��M�M��UR�EP�M�Q�p3�B���  �у���UR�EP��������]��������U����} w�E   �=p3 t$�EP�MQ�UR�p3�H���   �҃��E��j�EP�E������E��M��M��E���]���U����} w�E   �=p3 tT�} t$�EP�MQ�UR�p3�H���   �҃��E��"�EP�MQ�UR�p3�H���  �҃��E��E��E��j�MQ�������E��E���]���������U��EP�p3�Q��Ѓ�]��������U��EP�p3�Q��Ѓ�]��������U��EP�p3�Q��Ѓ�]��������U��EP�p3�Q��Ѓ�]��������U����  ��4����} u3��4����M���P�Q�P�Q�P�Q�P�Q�@�A�E��  �MQ��4���R�E�P��  ����4����QP��0�����0�����  ��0����$�lM j j �M���A�$�U����$�EP��4�����Q�U�R��  ��P�EP��4���Q�U�R�N  ��P��p���P�M�KM ��M�P�U�H�M��P�U�H�M��P�U���  �E�P�M���A�$�U����$�EP��4�����Q��X���R�>  ��P�EP��4���Q��@���R��  ��P��(���P�M�@M ��M�P�U�H�M��P�U�H�M��P�U��}� ��  �����$�����$�����$������ ���P�EP��4���Q������R�H  ��P������P�M�  P�MQ��4�����R��4���P������Q��  ��P������R�  ��P������P�M�p  P������Q��  ��P��h���R�s  ��P�E�P�  ���MQ��4���R��P���P�  ��P�M�Q�UR��4���P��8���Q�  ��P�� ���R�M��  P�����P�-  ��P������Q�M�:  P������R�]  ��P������P��  ����MȋP�ŰH�MЋP�UԋH�M؋P�U�j j �E���@�$�M����$�U�R�EP��4���Q������R��  ��P������P�M��J ��M�P�U�H�M��P�U�H�M��P�U��  �E�@��������D{8�MQ��x���R�M�b  ��M�P�U�H�M��P�U�H�M��P�U��q�E�P��H���Q�M�  ���@�$�U���B�$�E��� �$��`��������P��0���Q�M��  ��U�H�M�P�U��H�M�P�U��@�E���  j �M���A�$�U����$�EP��4�����Q�����R�  ��P�EP��4�����0Q�� ���R�  ��P������P�M�J ��M�P�U�H�M��P�U�H�M��P�U���4�����0P�M�Q������R�V  ��P������P��	  ��P��4������AH�$������R�
  ��P��4�����0P������Q�
  ����U�H�M�P�U��H�M�P�U��@�E��  j�MQ��4�����0R��p���P�  ��P�M�H ��4����IH�]��E���������Dz	�P��]��UR��4�����0P��X���Q�m  ��P��@���R�M��  P�EP��(���Q�Y
  ����U�H�M�P�U��H�M�P�U��@�E����]����E��$�M�Q�L  ����$�A  ���]��U�R�����P�  ��P���E��$������Q�R	  ����U�H�M�P�U��H�M�P�U��@�E��E��u����$�  �$��  �����M��]��MQ��4�����0R������P�n
  ��P������Q�M��  P�U�R������P�
	  ��P������Q�M�  ��U�H�M�P�U��H�M�P�U��@�E��MQ��8���R�
  ��P�E�P�MQ��	  ���E��]� �I �F =G �I iJ ~K U��Q�M���]� ���U����   ��<����}t
�   �Q  �M��I����EP��<������<����Bx�ЉEă}� u
�   �  �MQ�M�  �E��M�(  �E�j/�U�R�** ��j�E�P�* ���M�Q�UR�M�I  �E�    �	�E����E��}���   �}� uj �M�Q�M��  �j �U�R�M��  �E�    �	�E���E�M�;M�}u�U�3�;U���;E�t�ݍ�@����R  ��@���Q�U�R�EP��<������<����B|�Ѓ}��u��@����  �j j��@���Q�M�  ��@�����  �z����5����   ��]� ����������U��Q�M��   ��]� ��������������U��Q�M���]� ���U��Q�M���]�$ ���U��Q�M�3���]� �U����   ��$���j�EP�,  ����t�����   �M�Q�M�K  �E������E�    �	�U����U��EP��$������$����Bx��9E���   ��@����  ��@���Q�U�R�EP��$������$����B|�Ѓ}��u��@�����  뗋MQ�UR�E�P��@���Q��(���R�#  ��P�M��  ��t%�E��E�j�MQ��+  ����u��@����  ���@����s  �3����E���]� �����U���<  �������M�)  P������P�M�9  P��H���Q�  ���M��1  j �M��  �������U�R�EP�MQ��������������P|�ҍE�P�MQ��H���R�EP������Q�M�� ������ԋ�
�H�J�H�J�H�J�H�J�@�B�MQ�UR����������������   ��ǅ����   �M��y  ��������]� �������������U��Q�M�3���]� �U��Q�M�3���]� �U��Q�M��   ��]�$ ��������������U��Q�M���]� ���U��Q�M���]� ���U��Q�M���]� ���U��Q�M�3���]� �U��Q�M�3���]� �U���   �M��  ��tj �EP�MQ�L�������u3��   j h   ������R�[�����j �EP�M Q�UR�EP������Q�z   ���E��c �U��t�E� d �E�� t�E��c �M��   t�E��c �U��t�E��c h   ������P�MQ�URj�V  ����]����������������U��EP�MQ�UR�EP�MQ�UR��������E�M���   �Uǂ�   �c �Eǀ�    d �Mǁ�   `c �Uǂ�   �c �Eǀ�   �c �Mǁ�   pc �Uǂ�   d �Eǀ�   �c ]��������U���E�]����Au�E��E]�������U����E�$�� ��]�����������U�����]����Az
�h��+��`��]����u�X�����E�$�a� ��]�������������U��E�M� �I�U�E�B�����$�M�U�A�
�E�M� �I����$�U�E�B�H�M�U�A�J����$�M艽���E]�����U��E�M� �	�U�E�B�H���M�U�A�J�����$�   ��]��������U����E�$�� ��]�����������U����E�M� �	�U�E�B�H���M�U�A�J�����$�������]��E���������Dz�����$�M�U   �E�?���u��]��E�@�M����$�M�A�M����$�U��M����$�M脼���E��]��������������U��Q�M��E��E��M��E�Y�U��E�Z�E���]� ������U��E�@�M���$�M�A�M���$�U��M���$�M�	����E]�����U��E�M�@�A���$�U�E�B�@���$�M�U�����$�M������E]�������������U��E�M�@�a���$�U�E�B�`���$�M�U��"���$�M�q����E]�������������U��E�M�@(�	�U�E�B@�H���M�U�AX�J�����$�E�M�@ �	�U�E�B8�H���M�U�AP�J�����$�E�M�@�	�U�E�B0�H���M�U�AH�J�����$�M�κ���E]����������U��E�M�@(�	�U�B�E�M�@@�I���U�E�BX�H�����$�M�U�A �
�E�@�M�U�A8�J���E�M�@P�I�����$�U�E�B��M��U�E�B0�H���M�U�AH�J�����$�M�����E]���������U���hVWj �M��^  �E�M�@8�IX�U�E�BP�H@��M�I�U�E�BP�H(�M�U�A �JX��E�H0���M�U�A �J@�E�M�@8�I(��U�JH���]��E���������Dz�M�  �E�s  ���u��]��E�M�@�IX�U�E�BP�H��M�I0�U�E�B�H8�M�U�A�J@��E�HH���M�U�AP�J@�E�M�@8�IX��U�
���M��]��E�M�@�I(�U�E�B �H��M�IH�U�E�B �HX�M�U�AP�J(��E����M�U�AP�J�E�M�@�IX��U�J���M��]��E�M�@8�I(�U�E�B �H@��M�	�U�E�B@�H�M�U�A8�J��E�H���M�U�A�J �E�M�@�I(��U�J0���M��]��E�M�@8�IX�U�E�BP�H@���M��]��M�U�AP�J(�E�M�@ �IX���M��]��U�E�B �H@�M�U�A8�J(���M��]��E�M�@@�IH�U�E�BX�H0���M��]ȋM�U�AX�J�E�M�@(�IH���M��]ЋU�E�B(�H0�M�U�A@�J���M��]؋E�M�@0�IP�U�E�BH�H8���M��]��M�U�AH�J �E�M�@�IP���M��]�U�E�B�H8�M�U�A0�J ���M��]�   �u��}�E_^��]�U���d�M��M��߶���M����Զ���M���0�ɶ���M���H辶�������$�����$�����$�M�讶���M����P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�M��i����M������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�M��!����M���0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�M��ٵ���M���H���P�Q�P�Q�P�Q�P�Q�@�A�E���]�����������U��Q�M��EP�M��=   �MQ�M����.   �UR�M���0�   �EP�M���H�   �E���]� �������U��Q�M��E���]� U����M�EP�M�Q�U�R�p3�Hh�Q,�҃��M���P�Q�P�Q�P�Q�P�Q�@�A�E��]� �������������U����M�EP�M�Q�U�R�p3�Hh�Q0�҃��M���P�Q�P�Q�P�Q�P�Q�@�A�E��]� �������������U����M�EP�M�Q�U�R�p3�Hh�Q8�҃��M���P�Q�P�Q�P�Q�P�Q�@�A�E��]� �������������U���L�M��M�������M���������M���0���������$�M��y����E��M��U�P�M��H�U�P�M��H�U��P�����$�M��C����E����MЉ�UԉP�M؉H�U܉P�M��H�U�P�����$�M��
����E���0�M���U��P�M��H�UĉP�MȉH�ỦP�E��p��XH�M��AP    �E���]�����U��Q�M���]������U��Q�M��EP�M�Q�p3�BH��   �у���]� �������U��Q�M��E�P�p3�Qd�B<�Ѓ���]�U��Q�M��EP�MQ�U�R�p3�Hd�Q�҃���]� �������U��Q�M��EP�MQ�U�R�p3�Hd�Qp�҃���]� �������U��Q�M��EP�MQ�UR�E�P�p3�Qd���   �Ѓ���]� ���������������U���dVW�M��E�P�p3�QH�M��B,�й   ���}�E_^��]� ���������U��Q�M��EP�MQ�UR�E�P�p3�Qd�B�Ѓ���]� ��U���`VWj �M������E�M�@�	�U��E�M�@0�I���U�E�BH�H���]��M�U�A �
�E�@�M�U�A8�J���E�M�@P�I���]��U�E�B(��M�A�U�E�B@�H���M�U�AX�J���]��E�M�@�I�U�E�B0�H ���M�U�AH�J(���]��E�M�@ �I�U�E�B8�H ���M�U�AP�J(���]��E�M�@(�I�U�E�B@�H ���M�U�AX�J(���]ȋE�M�@�I0�U�E�B0�H8���M�U�AH�J@���]ЋE�M�@ �I0�U�E�B8�H8���M�U�AP�J@���]؋E�M�@(�I0�U�E�B@�H8���M�U�AX�J@���]��E�M�@�IH�U�E�B0�HP���M�U�AH�JX���]�E�M�@ �IH�U�E�B8�HP���M�U�AP�JX���]��E�M�@(�IH�U�E�B@�HP���M�U�AX�JX���]��   �u��}�E_^��]�������U��Q�M��EP�M�Q�p3�B@�H8�у���]� ����������U��Q�M��p3�PH�M��B$�Ћ�]������U���dVW�M��E�P�p3�QH�M��B<�й   ���}�E_^��]� ���������U��Q�M��M��   ����؋�]��������U��Q�M��p3�P�M��B<�Ћ�]�����̋�`L����������̋�`\����������̋�`l����������̋�`P����������̋�``����������̋�`p����������̋�`D����������̋�`T����������̋�`d����������̋�`t����������̋�`H����������̋�`X����������̋�`h�����������U��p3�H���   ��]������������U��E�Q�p3�B���   �у��U�    ]���������U��Q�M��E�P�p3�Q���   �Ѓ���]��������������U��Q�M��EP�M�Q�p3�B���   �у���]� �������U��p3�H���]����������������U��E�Q�p3�B�H�у��U�    ]������������U��E�Q�p3�B�H�у��U�    ]������������U����M�h�  �E�P�M�Q�p3�B���   �у����  �E��M���  �E���]��������������U��Q�M��E�P�p3�Q�B�Ѓ���]�U��Q�M��EP�M�Q�p3�B�H\�у���]� ����������U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�H���   �҃���]� ��������U��Q�M��EP�MQ�UR�EP�M�Q�p3�B�HX�у���]� ��������������U��Q�M��E�P�p3�Q�B �Ѓ���]�U��Q�M��EP�MQ�UR�EP�M�Q�p3�B���   �у���]� �����������U��Q�M��EP�MQ�UR�E�P�p3�Q�B�Ѓ���]� ��U��EP�MQ�UR�EP�MQ�p3�B��   �у�]����U��Q�M��EP�MQ�UR�EP�p3�Q�M��B$�Ћ�]� ��U��Q�M��EP�MQ�p3�B�M���x  �ҋ�]� �������U��Q�M��p3�P�M���|  �Ћ�]���U��Q�M��EP�MQ�UR�EP�M�Q�p3�B�H(�у���]� ��������������U��Q�M��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P�p3�Q�B`�Ѓ�(��]�$ ����������U��Q�M��EP�MQ�UR�EP�M�Q�p3�B�H,�у���]� ��������������U��Q�M��EP�MQ�UR�M�������P�M��٪����Pj j �E�P�p3�Q�B4�Ѓ� ��]� ������U��Q�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�p3�B�H4�у� ��]� ��U��Q�M��EP�MQ�U�R�p3�H�Q@�҃���]� �������U��Q�M��EP�M�Q�p3�B�HD�у���]� ����������U��Q�M��E�P�p3�Q�BL�Ѓ���]�U��Q�M��E�P�p3�Q�BL�Ѓ���]�U��Q�M��E�P�p3�Q�BP�Ѓ���]�U��Q�M��EP�M�Q�p3�B�HT�у���]� ����������U��Q�M��EP�M�Q�p3�B�HT�у���]� ����������U��Q�M��EP�MQ�U�R�p3�H���   �҃���]� ����U����M�EP�MQ�U�R�E�P�p3�Q���   �Ѓ�P�M�:  �M���  �E��]� ���������U��Q�M��E�P�p3�Q�Bh�Ѓ���]�U���h��h�   h�3h�   ��������E��}� t�M��m   �E���E�    �E���]�����������U����E�8 t*�M��U��E��E��}� tj�M���  �E���E�    �M�    ��]������������U��Q�M��M�����  �M��6   �E���]����������������U��Q�M��M��a   �M�����  ��]���U��Q�M��E��     �M��A`    �U��Bd    �E��@h    �M����Yp�U��Bx�����E��@|   ��]���U��Q�M��E��8 t j j j�M���Q�U��
�  �E��     �M��y` t�U���`R��������]������U��Q�M��E�P�M���dQ�U��BxP�MQ�U���`R�w������M��A|�U��z|u�E��8 u>�M��9 u�U��z|u
�E��@|�����M��    �U���`R�������E��@|�   �M��yd ��   �U���pR�E���hP�MQ� ����u$�U��Bh    �E����Xph��h  �  ���MQ�M����Q�  j j j�U���R�E���j  �M��A|�U��z|t�M������E��@|��M��Ax�����U��B|��]� �����U��Q�M��M��q����M�������]������U��Q�M��E��xd u�M��A`�}�U��E;Bxu�M��A`�j�UR�E��H`Qj�U���R�E����  �M��A|�U��z|u �E��M�Hx�} t	�U�   �E��@`��M��Ax�����} t�U�E��H|�
3���]� �����U��Q�M��} t�E�M��Ap��U��zd t�E��@h��M��y|u�   �3���]� ���������������U��p3�H���]����������������U��E�Q�p3�B�H�у��U�    ]������������U��Q�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�p3�B�H�у� ��]� ��U��Q�M��EP�M�Q�p3�B�H�у���]� ����������U��Q�M��E�P�p3�Q�B�Ѓ���]�U��Q�M��EP�MQ�U�R�p3�H�Q�҃���]� �������U��QV�M��EP�MQ�UR�M��d������M��Z����H �F@��^��]� �����������U��QV�M��EP�MQ�UR�M��$������M������H �FD��^��]� �����������U��QV�M��M�������xH u3���M���������M�������H �FH��^��]��������U��QV�M��M������xL u3��&�EP�MQ�UR�M��������M������H �FL��^��]� ���������U��QV�M��M��`����xP u����*�EP�MQ�UR�EP�M��=������M��3����H �VP��^��]� ����U��QV�M��M������xT u����"�EP�MQ�M���������M�������H �VT��^��]� ������������U��QV�M��M�������xX u�����EP�M��������M������H �VX��^��]� U���,V�Mԃ} t3�M��x�  �E�P�M��l������M��b����H �VL�ҋM��M����  �} t9�M��/���P�M��	  �M��n����M��&����P@�U�}� t�E�P�M�	  ^��]� �������U��QV�M��M�������x` u� }  ��EP�M���������M�������H �V`��^��]� ��������������U��QV�M��EP�M��������M������H �VH��^��]� ���U���V�M�j�EP�K	  �������P�M��Y����E��M螠��;E��M豠��;E�~������*�MQ�UR�EP�MQ�M��������M������H �VD��^��]� ����U��QV�M��M�������xP u������2�EP�MQ�UR�EP�MQ�UR�M���������M������H �FP��^��]� ����������U��QV�M��M������xT u������"�EP�MQ�M��s������M��i����H �VT��^��]� ����������U��QV�M��M��@����xX u��EP�M��,������M��"����H �VX��^��]� ���U����M���  �E�P�MQ��  ����t�}� u3���U�R�E�P�M�Q�U�R�M��������]���������U����M��M�?  �M��'�����uh��h�  �  ��3��   �E�    �E�P�M�Q�UR�E�P�p3�Q���   �Ѓ���u3��M�E�    �	�M����M��U�;U�}"�E��M�<� u��U��E��Q�M�]  �͍U�R�������   ��]� ����U����M�M�  �M��g�����uh�h�  �T  ��3��   �E�    �E�P�M�Q�UR�E�P�p3�Q���   �Ѓ���u3��o�}� u3��e�E�    �	�M����M��U�;U�}:�E��M�<� t�U��E���������u�ϋM��U���E��M�Q�M�  뵍U�R��������   ��]� ��U��p3�H��   ��]������������U��E�Q�p3�B��$  �у��U�    ]���������U��Q�M��E�P�MQ�p3�B��(  �у��E���]� ����U��Q�M��E�P�MQ�p3�B��,  �у���]� �������U��Q�M��E�P�MQ�p3�B��,  �у��������]� U��p3�H��0  ��]������������U��p3�H��4  ��]������������U��p3�H��p  ��]������������U��p3�H��t  ��]������������U����M��} t�M�yk  �E���E�    �E�P�M�Q�p3�B��8  �у���]� �����������U��Q�M��EP�M�Q�p3�B��<  �у���]� �������U��Q�M��EP�MQ�UR�E�P�p3�Q��@  �Ѓ���]� ���������������U��Q�M��EP�MQ�U�R�p3�H��D  �҃���]� ����U��Q�M��EP�M�Q�p3�B��H  �у���]� �������U����M�EP�M�Q�U�R�p3�H��L  �҃�P�M�����M�觗���E��]� ��������������U��Q�M��E�P�p3�Q��T  �Ѓ���]��������������U��Q�M��EP�M�Q�p3�B��l  �у���]� �������U��Q�M��E�P�p3�Q��P  �Ѓ���]��������������U��Q�M��EP�M�Q�p3�B��X  �у���]� �������U��p3�H��\  ��]������������U��E�Q�p3�B��`  �у��U�    ]���������U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�H��d  �҃���]� ��������U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�H��h  �҃���]� ��������U��Q�M��E�P�p3���   ��Ѓ���]���������������U��Q�M��E�P�p3���   �B8�Ѓ���]��������������U��Q�M��E��     �M��A    j �UR�E�P�p3���   �B�Ѓ��E���]� ���������������U��Q�M��M��q����E��t�M�Q�������E���]� ����U����M��M��r  �E�    �	�E����E��}�}�M��U��D�    ��E���]�U��Q�M��M��s  ��]��������������U��EP�MQ�p3�B��0  �у�]����������������U��Q�M��E�P�MQ�p3�B�H�у��E���]� �������U��E#E]������U��Q�M��E��     �M��A    �U��B    �E��@    �M��A    �U��B    �E���]��������U����M�j�M��-  �E��EP�M�Q�  ���E�3�t�E�H���U�J�E���]� �����������U����M��E��8 t�M��Q���U��	�E����E��}� |��M��A    ��]���U����M�j�M��   Pj�E   ���E��}� t�EP�  ���M����E��E���E�    �E��]� ��������������U��E]���������U����EEk��+����E��E���}�U��}� u�}� u�E+E�E��E��E���]�U����M�E�HM�M��U�B�M����E��M�U�;Q��   j�EP�M�QR�y������E�E�P�M���Q�U�P�M���   P�  ���E��}� tW�M��u-�U�: t%�E�HQ�U�R�E�Q�2  ���U�R�  ���E�M���U�E�B�M�Q�E����M��	�U�B�E��M�U��Q�E���]� ������U����EPj�������E��}� t�M��U���M��M���E�    �E���]����U��Q�M��E���]���U��Q�M��E��M��U��E�B�E���]� ���������������U��M�e: P�M�,   P�EP�MQ�p3�B��  �у�]��������������U��Q�M��E��@%��� ��]�����������U��E��P�MQ�UR�ـ ��]�����U����E� h�   h@��M��2���P�MQ�UR�T�������]��������������U��E]���������U��Q�E��M��U�R軿�����E�     ��]������������U����M�M�b  �E��}�NIVbP�}�NIVb��   �}�TCAb,�}�TCAb�7  �}�$'  �j  �}�MicM��   �p  �}�INIbtJ�b  �}�atni$�}�atnit)�}�ckhc�  �}�ytsdtL�5  �}�cnyst�'  ��  �  �E�x t
�   �  �M��A   �U��M�P����   �E��M�B�ЋM��A    ��   �U�z u
�   ��   �E��M�B���   j hIicM�M�����E��MQ�U�R�E��M�B���   j hIicM�M�S����E��MQ�U�R�E��M�B���Zj hdiem�M�*����E��MQ�U�R�E��M�B�ЉE��E��+�M��M�B�����MQ�U��M�P�Ҹ   �3���]� ���������U��Q�M��E�� ���M�QhP� �p3�B0��у��U��B�E��@    �E���]�U���,�E�    �M����  �} tO�EP�p3�Q4�B�Ѓ��E�}� u�E�    �M��8�  �E��   �M�Q�UR�E��M�B(�ЉE��J�MQ�p3�B0�H�у��E��}� u�E�    �M����  �E��N�U�R�EP�M���M��B �ЉE��M��_  ���t�M�Q�UR�p3�H0�Qx�҃��E��EԍM���  �Eԋ�]���U��Q�M��E�� ���M��y t�U��BP�p3�Q0�B�Ѓ��M��A    ��]��U��Q�M��E��HQ�p3�B0���   �у���]�����������U��Q�M��EP�M��QR�p3�H0���   �҃���]� �����U��Q�M��M��!_  P�p3�H0���   �҃���]����������U��Q�M�j j j j j j j j j4�E��HQ�p3�B0���   �у�(��]���������U��Q�M�j j j j j j j j j;�E��HQ�p3�B0���   �у�(��]���������U��Q�M��EP�M��m^  P�p3�Q0���   �Ѓ���]� ��U��� �M��E P�M����  �MQh8kds�M��Z����E�    �U�R�E�Pj �MQ�UR�EP�MQ�URj2�M���]  P�p3�H0���   �҃�(�E��E�M���  �E��]� U��Q�M��M���]  P�p3�H0���   �҃���]����������U��Q�M��E��x u3��aj j j j j �M Qj �URj�E��HQ�p3�B0���   �у�(�UR�EP�MQ�URj �EP�M��QR�p3�H0���   �҃���]� �����U��Q�M��E��x u3���M��QR�p3�H0�Q�҃���]��U��Q�M��M��������]� �����������U����M�E�x uj �M�]  �E�I�M�\  P�MQ�M�*3 P�U�BP�M�Q�p3�B0���   �у�P�M�A����M�������E��]� U��Q�M��EP�M��QR�p3�H0�Q�҃���]� ��������U��Q�M��E��x u�/j j j j j j �MQj j�U��BP�p3�Q0���   �Ѓ�(��]� ���������U��Q�M��E��x u3��.�M��[  P�MQ�M�G2 P�U��BP�p3�Q0�B�Ѓ���]� ��������U��Q�M��E��x u3��,�M�t[  P�M��1 P�M��QR�p3�H0���   �҃���]� ����������U��Q�M��E��x u3��.�M�$[  P�MQ�M�1 P�U��BP�p3�Q0�B\�Ѓ���]� ��������U��Q�M��E��x u3��#�MQ�UR�E��HQ�p3�B4��  �у���]� ���U��Q�M��E��x u3�� �MQ�UR�E��HQ�p3�B4�Hh�у���]� ������U��Q�M��E��x u3�� �MQ�UR�E��HQ�p3�B4�Hp�у���]� ������U��Q�M��E��x u3��#�MQ�UR�E��HQ�p3�B4��  �у���]� ���U��Q�M�h���h  ��EPj 3Ƀ} ����Qj �UR�EP�M��
   ��]� ����U���,�M�htniv�M����  �EPhulav�M�蹉��hgnlfhtmrf�M�觉���MQhinim�M�薉���URhixam�M�腉���EPhpets�M��t����MQhsirt�M��c����}   �u	�}$���t"�U Rh2nim�M��@����E$Ph2xam�M��/����M�Q�UR�E�P�M������������E�M��I����M���  �E��]�  ��������U���,�M�htlfv�M��
�  ���E�$hulav�M��X  �E,Phtmrf�M�賈�����E�$hinim�M��X  ���E�$hixam�M��wX  ���E$�$hpets�M��aX  �MDQhsirt�M��`����E0��������Dz�E8��������D{,���E0�$h2nim�M��X  ���E8�$h2xam�M��X  �U@Rhdauq�M������E�P�MQ�U�R�M���������\����E�M��!����M��i�  �E��]�@ U���T�M�hgnrs�M����  �EP�M���W  �M�Qj�M���W  �M�������UR�M��W  �E�Pj�M���W  �M������M�Q�UR�E�P�M��b�����������EčM������M����  �Eċ�]� ���������������U���,�M�hmnrs�M��J�  �EPj�M������M�Q�UR�E�P�M���������a����E�M��&����M��n�  �E��]� �����U���,�MԋE�����DSSSP�M����  j�M��%V  P�M�蜆���M�Q�UR�E�P�M�������������E�M������M����  �E��]� �����U���,�M�hCITb�M��z�  �EPhCITb�M��Y����MQhsirt�M��(����URhulav�M������E�P�MQ�U�R�M��������l����E�M��1����M��y�  �E��]� U����M�j �EP�M�Q�M�b  P�UR�M��X����E��M������E���]� ����U��Q�M��E,Pj �����$�����$htemf���E$�$���E�$���E�$���E�$�MQ�M��^�����]�( ��������U����M��E���������Dz�E�]�����E�$�U  ���]��E���������Dz�E�]�����E�$�aU  ���]�E,Pj �����$�����$hrgdf���E$�$�2U  �$���E��$���E��$���E�$�MQ�M�������]�( ��U��Q�M��E,Pj �����$�����$htcpf�E$�5p����$�E�5p����$�E�5p����$���E�$�MQ�M��,�����]�( ������U��Q�M��E��x u3��D�M��S  P�M Q���E�$���E�$�UR�M�1* P�E��HQ�p3�B0�H(�у�$��]� ��U����M�E�x u3��B�M�bS  P�M�Q�M��) P�U�BP�p3�Q0�B,�Ѓ��E�3Ƀ}� ���U�
�E���]� ��U��Q�M��E��x u3��.�M�S  P�MQ�M�) P�U��BP�p3�Q0�B,�Ѓ���]� ��������U��Q�M��E��x u3��.�M�R  P�MQ�M�7) P�U��BP�p3�Q0�B0�Ѓ���]� ��������U��Q�M��EP�MQ�M�������u3��;�U��R�EP�M��~�����u3�� �M��Q�UR�M��c�����u3���   ��]� U����M�E�x u3��   �E�    �M��Q  P�M�Q�M�{( P�U�BP�p3�Q0�B8�Ѓ��E��}� tG�}� tA�M�Q�M�����}� t(�U��U��E��E�}� tj�M��eR  �E���E�    �E�    �E���]� ���������U��� �M��M������E�P�MQ�M��/����E��}� u�E�    �M��~���E���U�R�M�^  �E��E�M��~���E��]� ���������������U��Q�M��E��x u3��2�M��P  P�MQ�UR�M�c' P�E��HQ�p3�B0�H<�у���]� ����U����M��E�    �E�P�MQ�M������E��U�R�EP�M�}Q  �E���]� ����U����M�E�P�MQ�M��7����E��U�R�EP�M�t����E���]� �����������U����M�E�P�MQ�M��G����E����E��$�UR�M�P  �E���]� ������U����M�M���~���E�P�MQ�M��������u3��E�U�R�EP�M��������u3��-�M�Q�UR�M��������u3���E�P�MQ�M�����   ��]� ������������U����M�M��~���E�P�MQ�M��/����E��U�R�EP�M����M��M�M��|���E��]� �����U���(�M؍M��Z  �E�P�MQ�M������E��U�R�EP�M�P  �M��M܍M���Z  �E܋�]� �����U���,�MԍM��}���E�P�M�Q�UR�M������E��}�t�E�P�MQ�M��~���}�t���E��$�UR�M�N  �E���]� ��������������U��Q�M�j j �EP�M�O  P�MQ�M��L�����]� ������U��Q�M��E$P�M Qj �UR�EP�MQj �UR�M��}��P�EP�M��H�����]�  ��U��Q�M�j �E@P���E8�$���E0�$�M,Q���E$�$���E�$���E�$�����$�UR�M�.O  ���$�EP�M��������]�< ������U��Q�M�j ���E$�$���E�$���E�$�����$�EP�M��N  ���$�MQ�M��������]�$ U��Q�M�j ���E$�$���E�$���E�$�����$�EP�M�N  ���$�MQ�M��������]�$ U��Q�M�j ���E$�$���E�$���E�$�����$�EP�M�8N  ���$�MQ�M��F�����]�$ U���(�M؋EPj �M��{��P�MQ�U�R�M�ؔ��P�EP�M��+����E��M���y���M��y���E���]� ���������������U���@�M�j �M��W  P�EP�M�Q�M��M  P�UR�M��O����E��M��X  �M��X  �E���]� ���U���<�M����]��}�t�����$�EP�M�HM  �]��M Q���E�$���E��$�M��z��P�UR�E�P�M�f{��P�MQ�M�������]� ���U���L�M̃} u�p3�H���   �҉E�} u3��y  �M�	 �E�htlfv�M���  �M�QM  �M���$�#M  ���M�]��EM  ���$�
M  ���}ă��$hulav�M��K  hmrffhtmrf�M���z���M��L  �M���$��L  ���M�]���L  ���$�L  ���}����$hinim�M��J  �M�L  �M���$�L  ���M�]��L  ���$�hL  ���}����$hixam�M��_J  �����$hpets�M��JJ  j hdauq�M��Kz���E�Phspff�M��:z���M Qhsirt�M��)z���U�R�EP�M�Q�M��������~����E�M��C����M���  �E��]� ��U���,�Mԃ} u�p3�H���   �҉E�} u3��`�M�l �E�E�P�MQ�M������E��E������$�E������$�M��p  �U��
�H�J�H�J�@�B�E���]� ��������������U���$�M�j �E P�MQ�UR�M��aK  P�EP�M�Q�M�pK  P�UR�EP�M��o�����]� ���������U����M�M��K  �E�P�MQ�UR�M�������E��E�P�MQ�M�hK  �E���]� ���������������U��Q�M��E��x u3��:�M�dH  Pj j j j j j �M�� Pj1�M��QR�p3�H0���   �҃�(��]� ������������U����M��E��x u3��B�E�    �M�Qj j �UR�EP�MQ�UR�EPj�M��QR�p3�H0���   �҃�(�E���]� ��U��Q�M��E��x u3��/j j j j j j j �MQj-�U��BP�p3�Q0���   �Ѓ�(��]� �������U����M��E��x u3��<�E�    �M�Qj j j �UR�EPj j j)�M��QR�p3�H0���   �҃�(�E���]� ��������U����M��E��x u3��<�E�    �M�Qj j �URj �EPj j j)�M��QR�p3�H0���   �҃�(�E���]� ��������U��Q�M��E��x u3��5j j j �MQ�UR�EPj �MQj/�U��BP�p3�Q0���   �Ѓ�(��]� �U����M��E��x u3��B�E�    �M�Qj j �UR�EP�MQ�UR�EPj'�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��B�E�    �M�Qj j �UR�EP�MQ�UR�EPj,�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��B�E�    �M�Qj j �UR�EP�MQ�UR�EPj�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��E�E�    �M�Qj �UR�EP�MQ�UR�EP�MQj�U��BP�p3�Q0���   �Ѓ�(�E���]� ���������������U��Q�M�j j j �EP�MQ�URj �EPj.�M��QR�p3�H0���   �҃�(��]� ���������������U����M��E��x u3��B�E�    �M�Qj �UR�EP�MQ�URj �EPj�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��B�E�    �M�Qj �UR�EP�MQ�URj �EPj:�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��B�E�    �M�Qj �UR�EP�MQ�URj �EPj�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��B�E�    �M�Qj �UR�EP�MQ�URj �EPj*�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��A�E�    �M�Qj j �UR�EP�MQj �URj�E��HQ�p3�B0���   �у�(�E���]� ���U����M��E��x u3��A�E�    �M�Qj j �UR�EP�MQj �URj�E��HQ�p3�B0���   �у�(�E���]� ���U����M��E��x u3��A�E�    �M�Qj j �UR�EP�MQj �URj	�E��HQ�p3�B0���   �у�(�E���]� ���U����M��E��x u3��A�E�    �M�Qj j �UR�EP�MQj �URj
�E��HQ�p3�B0���   �у�(�E���]� ���U����M��E��x u3��B�E�    �M�Qj �UR�EP�MQ�URj �EPj�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��B�E�    �M�Qj �UR�EP�MQ�URj �EPj�M��QR�p3�H0���   �҃�(�E���]� ��U��Q�M��E��x u3��5j j j �MQ�UR�EPj �MQj�U��BP�p3�Q0���   �Ѓ�(��]� �U����M��E��x u3��B�E�    �M�Qj �UR�EP�MQ�URj �EPj�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��B�E�    �M�Qj �UR�EP�MQ�URj �EPj>�M��QR�p3�H0���   �҃�(�E���]� ��U����M��E��x u3��A�E�    �M�Qj j �UR�EP�MQj �URj�E��HQ�p3�B0���   �у�(�E���]� ���U��Q�M��E��x u3��?�M�4?  Pj j j j �MQ�UR�M� Pj�E��HQ�p3�B0���   �у�(��]� �������U����M�EP�M����  �M�Q�U�R�M��K�  ��t+�}� u��M��w���P�E�P�MQ�M��V�����u3�����   ��]� �U��Q�M��E��x u3��:�M�t>  Pj j j j j j �M�� Pj�M��QR�p3�H0���   �҃�(��]� ������������U����M��E��x u3��A�E�    �M�Qj j �UR�EP�MQj �URj�E��HQ�p3�B0���   �у�(�E���]� ���U��Q�M��E��x u3��#�MQ�UR�EP�M��QR�p3�H0�QD�҃���]� ���U��Q�M��E��x u3��;�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E��HQ�p3�B0���   �у�$��]�  �����������U��Q�M��E��x u3���M��QR�p3�H0�QX�҃���]��U��Q�M��E��x u3�� �MQ�UR�E��HQ�p3�B0�HL�у���]� ������U��Q�M��E��x u3��"�M��   �Q�U��BP�p3�Q0�BP�Ѓ���]� ����U��Q�M��E��x u3���MQ�U��BP�p3�Q0�BP�Ѓ���]� ����������U��Q�M��E��x u3��(�MQ�UR�EP�MQ�U��BP�p3�Q0�BT�Ѓ���]� ��������������U��Q�M��E�HQ�p3�B4��у��U�B    �E�M��H�M�;  P�UR�EP�M�6 P�M��QR�p3�H0���   �҃��M�A�U3��z ����]� ���U��Q�M��E��x u3��/j j j j j �MQj j j�U��BP�p3�Q0���   �Ѓ�(��]� �������U��Q�M��} u3��4�E�@    �M��:  P�MQ�M���:  P�p3�B0���   �у���]� �����U��Q�M�j j j j j j j j j0�M��:  P�p3�H0���   �҃�(��]��������U��Q�M��} u�E`3�EP�M�  P�MQ�U��BP�p3�Q0�B@�Ѓ���]� �������������U��Q�M��EP�MQ�UR�EP�MQ�U��BP�p3�Q0�Bd�Ѓ���]� �������U��Q�M��EP�MQ�UR�EP�MQ�U��BP�p3�Q0�Bp�Ѓ���]� �������U��Q�M��M�9  P�EP�MQ�UR�EP�M�( P�M��QR�p3�H0�Qh�҃���]� ����������U��Q�M�j j j j j j j �M�� Pj�E��HQ�p3�B0���   �у�(��]� ���������������U��Q�M�j j j j j jj �M� Pj�E��HQ�p3�B0���   �у�(��]� ���������������U��Q�M�j j j j j j j �M�C Pj�E��HQ�p3�B0���   �у�(��]� ���������������U��� �M��M�蟾  �M�g8  P�E�Pj j j j j �M�� Pj8�M��QR�p3�H0���   �҃�(�E�}� t�E�P�M���  �M�M�M��о  �E��]� �������U��Q�M��M��7  P�EPj j j j j �M�j Pj9�M��QR�p3�H0���   �҃�(��]� �������U��Q�M��M�7  Pj j j j j j �M� Pj"�E��HQ�p3�B0���   �у�(��]� ��������U��Q�M��M�Q7  Pj j j j j j �M�� Pj5�E��HQ�p3�B0���   �у�(��]� ��������U��Q�M��M�7  Pj j j j �EPj �M�z Pj<�M��QR�p3�H0���   �҃�(��]� �������U��Q�M�j j �EP�MQ�UR�EPj �MQj3�U��BP�p3�Q0���   �Ѓ�(��]� ������������U��Q�M�j j j j j �EPj �MQj�U��BP�p3�Q0���   �Ѓ�(�MQ�U��BP�p3�Q0�Bt�Ѓ���]� ������U��Q�M�j j j j j j �EPj j�M��QR�p3�H0���   �҃�(��]� �����U��Q�M�j j j j j j j j j�E��HQ�p3�B0���   �у�(��]���������U��Q�M�j j j j j j j �EPj�M��QR�p3�H0���   �҃�(��]� �����U��Q�M�j j j j j j j j j(�E��HQ�p3�B0���   �у�(��]���������U��Q�M�j j j j j j �EP�MQj&�U��BP�p3�Q0���   �Ѓ�(��]� ��U��Q�M�j j j j �EP�MQj �URj+�E��HQ�p3�B0���   �у�(��]� U��Q�M�j j j j j j j j j�E��HQ�p3�B0���   �у�(��]���������U��Q�M�j j j j j j j j j#�E��HQ�p3�B0���   �у�(��]���������U��Q�M��} tj j�M��c���M��} tj j�M�c���U��EP�MQ�U��BP�p3�Q0�B`�Ѓ���]� �����U��Q�M��EP�MQ�UR�E��HQ�p3�B0���   �у���]� ������������U��Q�M�j j j j j j j j j �E��HQ�p3�B0���   �у�(��]���������U��Q�M��   ��]�U��Q�M��   ��]�U��Q�M���]������U��Q�M��   ��]� ��������������U��Q�M�3���]� �U��Q�M�3���]����U��Q�M���]� ���U��Q�M��M������E�� ��M��A   �U��B    �E���]��������������U��Q�M��E�� ��M�������]�����U����M��E��@    j �MQ�UR�EP�MQj 3҃} ��
R�M��t�����t�E��x t	�E�   ��E�    �E���]� ��������������U��Q�M��E��M�H�M�������]� ��U����M�M�_1  �E��}�ckhc �}�ckhct,�}�cksatS�}�TCAbtf��   �}�atnit�   3��   �E�x t �M��������t�M��A    �   �   3��   �U�z t�E��M�B���t3��pj hdiem�M��`���E��M��A   �UR�E�P�M��M�B�ЉE��M�y t�}�t�}�u3҃}���R�M�������E���EP�MQ�M��������]� ������������U����M�E�x u��   �M�M��}���   �U��$��� �E;E~��   �   �M;M|�   �{�U;U}�   �l�E;E�   �]�M;M~�U;U}�   �F�E;E|
�M;M�v�2�U;U|
�E;E}�b��M;M~
�U;U�N�
�E;Et�B�MQ�M���2  �U�R�M������j�E���$�E���$�EP�>�  ���M��A    ��]� �I �� �� ² Ѳ � �� � � 3� ����U����M�E�x u�I  �M�M��}���   �U��$�� �E�]����z�  ��   �E�]����Az�  �   �E�]����Au��   �   �E�]����u��   �   �E�]����z�E �]����Au�   �n�E�]����Az�E �]����u�   �M�E�]����Az�E �]����Au�u�/�E�]����z�E �]����u�W��E�E������D{�D�EP�M��h1  �M�Q�M��\����U(R���E �$���E�$�EP��  ���M��A    ��]�$ ��� �� � &� =� ^� � �� �� ����U��Q�M�j���E �$���E�$���E�$�EP�MQ�M��<�����]�  ������U��Q�M�j���E �$���E�$���E�$�EP�MQ�M��������]�  ������U��Q�M�j���E �$���E�$���E�$�EP�MQ�M�������]�  ������U��Q�M��E�� D��M��A    �U��B    �E��@    �E���]������������U��Q�M��E�� D��M��y u�U��BP�p3�Q4��Ѓ��M��A    �U��B    ��]���������U��Q�M��EP�M��QR�p3�H4�Qt�҃���]� ��������U����M��} tA�EP�M��5,  P�p3�Q0���   �Ѓ��E��MQ�U�R�p3�H0���   �҃���EP�M��QR�p3�H0�Q|�҃���]� ���������������U��Q�M��E��HQ�p3�B4�H�у���]��������������U��Q�M��E��HQ�p3�B4�H�у���]��������������U��Q�M��E��HQ�p3�B4�H�у���]��������������U��Q�M��E��HQ�p3�B4�H|�у���]��������������U��Q�M��E��HQ�p3�B4���   �у���]�����������U��Q�M��E$P�M Q�UR�EP���E�$���E�$�M��QR�p3�H4��  �҃�$��]�  �������U��Q�M��EP�MQ�UR�EP�M��QR�p3�H4�Q�҃���]� ������������U��Q�M��EP�MQ�UR�EP�M��QR�p3�H4�Q�҃���]� ������������U��Q�M��M�-  ��u�M�-  P�M��;   �2�M�q-  ��u�M�t���P�M��K   �h��h
  �j�������]� �U��Q�M��EP�M��QR�p3�H4�Q �҃���]� ��������U��Q�M��EP�M��QR�p3�H4�Q$�҃���]� ��������U��Q�M��EP�MQ�UR�EP�M��QR�p3�H0���   �҃���]� ���������U��Q�M��EP�M��QR�p3�H0���   �҃���]� �����U��Q�M����E�$�EP�MQ�U��BP�p3�Q0���   �Ѓ���]� �������U��Q�M��EP�M��QR�p3�H4���   �҃���]� �����U��Q�M��EP�MQ�UR�EP�MQ�U��BP�p3�Q4���   �Ѓ���]� ����U��Q�M��EP�MQ�UR�EP�MQ�U��BP�p3�Q4���   �Ѓ���]� ����U��Q�M��EP�M��QR�p3�H4�Q(�҃���]� ��������U��Q�M��EP�MQ�UR�E��HQ�p3�B4�H,�у���]� ���������������U��Q�M��EP�MQ�U��BP�p3�Q4�B0�Ѓ���]� ���U��Q�M��E��HQ�p3�B4�H4�у���]��������������U���0�M��E�    �E�    �E�P�M�Q�UR�E܋H������M��z���P�M��*  �M�Q�U�R�E�P�M�Q�U�R�E܋H�����} tC�} t=�M�;M�~'�U�U�9U�}�E�;E�~�M�M�9M�}	�E�   ��E�    �E��V�.�} t(�U�;U�~�E�E�9E�}	�E�   ��E�    �E��&�M�;M�~�U�U�9U�}	�E�   ��E�    �EЋ�]� ���������������U��Q�M��EP�M��QR�p3�H4�Q8�҃���]� ��������U��Q�M��EP�M��QR�p3�H4�Q<�҃���]� ��������U��Q�M��EP�MQ�U��BP�p3�Q4���   �Ѓ���]� U��Q�M����E�$�E��HQ�p3�B4��  �у���]� ���������������U��Q�M��E��HQ�p3�B4�H@�у���]��������������U��Q�M��E��HQ�p3�B4��  �у���]�����������U��Q�M��EP�MQ�U��BP�p3�Q4�BD�Ѓ���]� ���U��Q�M��EP�MQ�U��BP�p3�Q4�BH�Ѓ���]� ���U��Q�M��EP�MQ�U��BP�p3�Q4�BL�Ѓ���]� ���U��Q�M��EP�MQ�U��BP�p3�Q4�BP�Ѓ���]� ���U��Q�M��M�'  ����   �M�'  ��u,�M�'  P�M�'  P�E��HQ�p3�B4�HP�у��K�M�W'  ��u,�M�Z���P�M�q'  P�U��BP�p3�Q4�BH�Ѓ��h��h�  �7������   �M�'  ����   �M��&  ��u+�M�'  P�M����P�M��QR�p3�H4�QL�҃��K�M�&  ��u,�M�����P�M踺��P�E��HQ�p3�B4�HD�у��h�h�  螻�����h(�h�  芻������]� �U��Q�M��EP�MQ�UR�EP�M��QR�p3�H4��  �҃���]� ���������U��Q�M��E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP�M��QR�p3�H4�QT�҃�,��]�( ����U��Q�M��EP�MQ�UR�EP�M��QR�p3�H4�QX�҃���]� ������������U��Q�M��E��HQ�p3�B4�H`�у���]��������������U��Q�M��E��HQ�p3�B4�Hd�у���]��������������U��Q�M��EP�MQ�UR�EP�M��QR�p3�H4��   �҃���]� ���������U��Q�M��EP�MQ�UR�EP�MQ�UR�E��HQ�p3�B4�H\�у���]� ���U��Q�M��EP�MQ�U��BP�p3�Q4�Bh�Ѓ���]� ���U��Q�M��EP�MQ�U��BP�p3�Q4��  �Ѓ���]� U��Q�M��EP�MQ�U��BP�p3�Q4��  �Ѓ���]� U��Q�M��EP�MQ�U��BP�p3�Q4�Bp�Ѓ���]� ���U���4�M̋Ẽx tp�} t(�M������P�M̋I�4   P�p3�B0�Hl�у��B�M�����P�M��?#  hARDb�M��b�  P�U�R�E�P�M̋I�����M��V����M�螦  ��]� ��������U��Q�M��EP�M��QR�p3�H4�Ql�҃��   ��]� ���U��Q�M��EP���E�$���E�$�MQ�U��BP�p3�Q4���   �Ѓ���]� ��������������U��Q�M��EP�MQ�UR�E��HQ�p3�B4���   �у���]� ������������U��Q�M��E��HQ�p3�B4���   �у���]�����������U��Q�M��E��HQ�p3�B4��  �у���]�����������U��Q�M��   ��]�U��Q�M��   ��]�U��Q�M�h�  �M�������EP�MQ�UR�EP�M�����2���]� ������������U��Q�M��EP�MQ�UR�EP�M���M��B�Ћ�]� ������U��Q�M��   ��]� ��������������U��Q�M�3���]� �U��Q�M���]� ���U��Q�M�3���]� �U��Q�M���]� ���U��Q�M��EP�MQ�UR�EP�M��QR�p3�H4�Qx�҃���]� ������������U��Q�M��EP�MQ�UR�E��H������]� ������������U��Q�M��} tj j�M�M���M��} tj j�M��L���U��EP�MQ�U��BP�p3�Q4�Bp�Ѓ���]� �����U���(�M��E�    �M�  �E؁}�INIbT�}�INIb��   �}�SACb,�}�SACb��   �}�$'  ��  �}�MicM��  ��  �}�ARDb��   �  �}�NIVb(�}�NIVbtJ�}�NPIb�:  �}�ISIb��   �~  �}�cnys�H  �l  �E܋�M܋B���E�   �S  �M܋�M܋B���E�   �:  �E�    �E�    �M�Q�U�R�E܋�M܋B�Ѕ�t �M�Q�U�R�E܋HQ�p3�B4�H�у��E�   ��   �M�����P�M������P�U܋�M܋P���E�   �   j j�M�IK���E�j j�M�:K���E�j j�M�+K���E�j j�M�K���E�EP�M�Q�U�R�E�P�M�Q�U܋�M܋P���E�   �V�EP�M܋�M܋B���F�MQ�U܋�M܋P$���E�   �)j hIicM�M�J���E��EP�M�Q�U܋�M܋P ����E���]� U��Q�M�h����h����h�����EP�MQh����h����h����h�����UR�M��������]� ������������U����M�hYALf�M�躠  P�M������M��	�  ��]������U��Q�M��M��1����E�� t��M��A   �E���]��������U��Q�M��E�� t��M��(�����]�����U����M��M�  �E��}�cksat6�}�ckhct�G�E��@   �M��F�����t�M��A    �   �03��,�U��z t�E���M��B���3���MQ�UR�M�葶����]� �����������U��EP�MQ�UR�EP�MQ�UR�p3�H���  �҃�]�U��EP�p3�Q0���   �Ѓ�]����U����EP�MQ�U�R�p3�H0���   �҃�P�M�"H���M��JF���E��]����U���<�M���G���E�    �	�E����E��   ����   j �U�k�
R�M�bH���E�j �E�k�
��P�M�KH���E�}� u�S�}� ~#j hH��M��E���M�Q�M��o  �M��E���U�R�E�P�M�Q�&�����P�M��J  �M��E���d����U�R�M�QG���M��yE���E��]���U��EP�MQ�p3�B0���   �у�]����������������U��EP�MQ�UR�EP�MQ�UR�p3�H0���   �҃�]�U��EP�p3�Q0���   �Ѓ�]����U��j0j ��  ��P�EP��  ��]���U��j0j �  ��P�EP�U����P�ޥ  ��]����������U���j0j �q  ��P�EP�MQ�U�R�U����P裥  ���M��hD����]�����U���j0j �1  ��P�EP�MQ�UR�E�P��U����P�_�  ���M��$D����]�U��j j��  ��P�EP�7�  ��3Ƀ�����]���������U��j j��  ��P�EP��T����P���  ��3Ƀ�����]����������������U���j j�  ��P�EP�MQ�U�R�T����P賤  ��3Ƀ����M��M��mC���E���]�������U���j j�1  ��P�EP�MQ�UR�E�P��T����P�_�  ��3Ƀ����M��M��C���E���]���U��EP�MQj �p3�B���   �у�]��������������U��EP�MQ�URj �p3�H���   �҃�]�����������U��Q�M��EP�MQ�UR�E��HQ�p3�B4�H,�у���]� ���������������U��Q�M��EP�MQ�U��BP�p3�Q4�B0�Ѓ���]� ���U��Q�M��E��HQ�p3�B4�H4�у���]��������������U����M�M�/  � �E��M�  �E��}� t�E�   �M�Q�U�R�EP�M��n�����]� ��������U��Q�M��E P�MQ�M��  P�UR�EP�MQ�M��  �R�EP�M��e�����]� ���������������U��Q�M��M�  P�E<P���E4�$���E,�$�M(Q���E �$���E�$���E�$�M�  ��� �$�UR�M��ߺ����]�8 ���������U��Q�M��M�  P���E �$���E�$���E�$�M�=  ��� �$�EP�M��ٽ����]�  ���U��Q�M��M��  P���E �$���E�$���E�$�M��  ��� �$�EP�M�������]�  ���U��Q�M��M�q  P���E �$���E�$���E�$�M�  ��� �$�EP�M��Y�����]�  ���U��Q�M��M�!  P�EP�MQ�UR�M�\  P�EP�MQ�M��������]� �����U��Q�M��EP�M��  P�M��  P�MQ�M�������]� �U��Q�M��E P���E�$���E�$�M��  P�MQ�M�������]� ��������U���(�M�E�P�M�Q�UR�M�������E�P�M�Q�U�R�E�P�MQ�M�������} tC�} t=�U�;U�~'�E�E�9E�}�M�;M�~�U�U�9U�}	�E�   ��E�    �E��V�.�} t(�E�;E�~�M�M�9M�}	�E�   ��E�    �E��&�U�;U�~�E�E�9E�}	�E�   ��E�    �E؋�]� ����U����M�E�E��}� u	�M���M�j hdiuM�M�@���E��}� u�   �G�U��E�;u3��9j hIicM�M�@��9E�uj h1icM�M�  ��t3���M��U���   ��]� ������U���hfnic�M�  �E��}� tj
�M��  ��t�Vhfnic�E�P�M�3  P�M��  �M���  �M��  ���t�M��  ��uhfnic�M�  �MQj
�M�N@����]�����������U��Q�M��EP�MQ�UR�EP�M���  P�p3�Q0���   �Ѓ���]� ������U��Q�M��M�  Pj j j �EP�MQj �M��  Pj=�U��BP�p3�Q0���   �Ѓ�(��]� ����U��Q�M��M�Q  P�EPj j j��MQj �M���  Pj=�U��BP�p3�Q0���   �Ѓ�(��]� ����U��Q�M�j j j j j j j j j6�M���  P�p3�H0���   �҃�(��]��������U����M�j �EP�M�  �E��M�Q�M��j  ��]� ����U����M�j �EP�M�Y>���E��M�Q�M��:  ��]� ����U����M�����$�EP�M��  �]����E��$�M���  ��]� ���������U���L�M��M��=���M��=��P�EP�M�Q�M��=����U�H�M�P�U��H�M�P�U��@�E����̋U��E�A�U��Q�E�A�U��Q�E��A�M��  ��]� �������������U���4�M̍M���  �M���  P�EP�M�Q�M��  ��U��H�M�P�U��@�E����̋U���E�A�U��Q�E��A�M��;  ��]� �����U���8�MȍM��?<���M��7<��P�EP�M�Q�M�vU��P�M��ݥ���M��e:���M��]:�����̍U�R�<���M���  �M��?:����]� ���������U����M��E;Eu&j htsem�M�p<����uj hrdem�M�]<����t3��<�E�    �MQ�M��  �U�R�E�P�M������u3���M�Q�M��  �   ��]� ���U����M��E;Eu&j htsem�M��;����uj hrdem�M��;����t3��<�E�    �MQ�M��"  �U�R�E�P�M�¸����u3���M�Q�M��  �   ��]� ���U����M�E;Eu&j htsem�M�p;����uj hrdem�M�];����t3��?���]��MQ�M��  �U�R�E�P�M蔸����u3�����E��$�M���  �   ��]� U���4�M̋E;Et�M;Mt�U;Ut3��   j htsem�M��:����uj hrdem�M��:����t3��   �����$�M��k}���EP�M���  �MQ�M���  �UR�M���  �E�P�M�Q�U�R�E�P�M������u3��5���̋U��E�A�U��Q�E�A�U��Q�E��A�M��g  �   ��]� ������������U����M�E;Eu&j htsem�M� :����uj hrdem�M��9����t3��Y�M��m  �MQ�M��1  �U�R�EP�M�Q�M�-�����u3��)���ԋE���M�J�E��B�M��J�M���  �   ��]� ������U���(�M؋E;Eu&j htsem�M�`9����uj hrdem�M�M9����t3��d�M��8���MQ�M��  �U�R�E�P�M�1�����u�E�    �M��6���E��(���̍U�R�k8���M��3  �E�   �M��6���E܋�]� �����������U��Q�M��M������E�� ���M��U�Qj hmyal�M�8���M��A�U��zt�E��xt
�M��A    j
hhfed�M�o8���U��B�E���]� U����M��M�/  �E��}�ytsdt��M�虪���E���M��B�и   ��MQ�UR�M��U�����]� ���������������U��Q�M�3���]����U��Q�M�3���]����U��Q�M���]������U��Q�M�3���]����U��Q�M�3���]����U��Q�M�3���]����U��Q�M�3���]� �U����M�M��  �E�P�M�s  �M��K  �E��]� ��U��Q�M��E���M��BD�Ѕ�t!�M��Q;Ut�E��M�H�U���M��PH�ҋ�]� �U��Q�M��E��@��]����������������U��Q�M��E��x u3���M��Q�������؋�]��������U��Q�M���]������U��Q�M��L���]�U��Q�M������$�E��H�6   �M�Q�U��B�M��I��B$��j j h���豘  ����]�����������U��Q�M��E��E�X(��]� ����������U���l�M��E�P�M���M��B(��P�M������M��3��j j j �M��W5��Pj jj?j �M������M��3��j �M��45��Pj j(�
  ��Pjh�  �M�����������EߍM��U3���M߅�t3��   j j j �M���4��Pj j j8j �M��'����M��3��j�M��%����M��͋  Pj�  ��Ph,  �  ��Pj;�M��4��Ph	��h�  �M������M���2���M���  �M������M�����j�M�������U��E��B$j��  ���   ��]�U����M�j�M���Z�  �E��@4    �M��A8    �U��B<    �E����X(h�   �M��w���j h\��M���1��h�  �M���  j j �M�Q�U�R�M��w����M��2��j j�M����  ��]�������������U��Q�M��E�����]����������������U����M��E�    �   ����   �M��y4 t4h`�h~  �ۜ����j
�1�  ���M����
  ��t3��   �ËM���0�+
  �U��z4 ur�E��M�H8�U��E�B4�M���0�%
  �M��y4 tj
�՞  ���M����'
  ��t3��T�؋M���0��	  �U��B<�E��M��A<    �M���0��	  �$�h��h�  �!������M���0�	  �����E���]� �����U���l�M�j h���M��h0��h�  �M��[  j j �E�P�M��A(�p�� P�U�R�x2����P�E�P�	  ��P�M�Q�M�軬���M��S0���M��K0���M��C0��htats�M��&�  jj�M��  �U����B(�$j�M���  h�  �M���  �E�P�M�Q�U�R�M�賥���M������E��x4 t_�M���0�  �M��y4 t.�U��B8P�M��Q4�҃��M��A<�U��B8    �E��@4    �h��h�  �њ�����M���0�c  �M��ˈ  ��]� �����U���L�M��M�  �E��}�MicMtq�}�ckhctD�}�fnict��   j�M��"�  P�M虈  �M��q�  jj�M��1���   �   �   �E���M��B�Ѕ�u3��   �   �   �qj hIicM�M�31���E��}����t�Thtats�M�訇  j j�M��<  h�  �M��_  �M�Q�U�R�E�P�M��K����M�胘���M��ˇ  j�M��!����MQ�UR�M��1�����]� �����������U����M��E�E��}�t�(j�M�����  j蕎  ��j �M�������   ��MQ�UR�M�������]� �����������U��Q�M�j�M�����  j�E�  ��3���]�������������U��Q�M��p3�P�M��B �Ћ�]������U��Q�M��M��Q����E��t�M�Q��_�����E���]� ����U��Q�M��E��@��]����������������U��Q�M����E�$�EP�p3�Q�M��B,�Ћ�]� �����U��Q�M��E��    �M��U�Q�E���]� ��������������U��Q�M��EP�MQ�p3�B�M����   �ҋ�]� �������U���E���5 �]�������������U��Q�M��M��,���E��t�M�Q��^�����E���]� ����U��Q�M��EP�MQ�p3�B�M��P0�ҋ�]� ����������U��Q�M��EP�MQ�p3�B�M��P<�ҋ�]� ����������U��Q�M��EP�MQ�p3�B�M����   �ҋ�]� �������U��Q�M����E�$�EP�p3�Q�M����   �Ћ�]� ��U��� �M��EP�MQ�U�R�p3�P�M����   ��P�M��	  �M��'
  �E��]� ��������������U����E�$� ��]�����������U��Q�M��E�� ��]�U��Q�M��E��@��]����������������U��Q�M��E�����M����Y�E���]����U����M�EP�MQ�U�R�p3�P�M싂�   �ЋM���P�Q�P�Q�@�A�E��]� ������U��Q�M��EP�MQ�p3�B�M��P@�ҋ�]� ����������U��Q�M��M������E��t�M�Q�\�����E���]� ����U��Q�M��E��M��U��B    �E���]� ��������������U��Q�M��M�������E��t�M�Q�P\�����E���]� ����U��Q�M��E�P�p3���   �B�Ѓ���]��������������U��Q�M��E�P�p3���   �B@�Ѓ���]��������������U��Q�M��M�������E��t�M�Q��[�����E���]� ����U��Q�M�j�j��EP�M���{��P�M��C���E���]� �������U��EE]������U��Q�M��EP�MQ�p3�B�M����   �ҋ�]� �������U��Q�M��EP�p3�Q�M��B$�Ћ�]� ��������������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U����M�EP�M�Q�p3�B�M�PP��P�M�u�  �M�蝁  �E��]� ����U��Q�M��EP�p3�Q�M��BT�Ћ�]� ��������������U��Q�M��M��!   �E��t�M�Q�PZ�����E���]� ����U��Q�M��M��Q�����]��������������U��Q�M��M���讑����]�����������U��Q�M��E��M���E��P�M����ݑ���E���]� ����U��j �EP�   ��]��������������U��E��E]���U��Q�M��p3�PP�M��Bh�Ћ�]������U��Q�M��p3�PP�M��Bl�Ћ�]������U��Q�M��E��HQ�p3�BP�H�у���]��������������U����EP�M��(���MQ�M��b����U�R�M�v(���M��&���E��]��������U����M�M���,   �E�� �����M��   P�M���?   �M��W����E��]�U��Q�M��E��     �M��A    �E���]����������������U��Q�M�j �E�P�M�   �E���]� ��U��Q�M��EP�M�Q�UR�p3���   �Q�҃���]� ����U��Q�M��E�����]����������������U��Q�M��E��8�u�M��    �U��E�B��M��9 u�U��B;Et	�M��   ��]� �����������U��Q�M��E��8�u�M��    �UR�M���詐���$�E��8 u�MQ�M����    ��t	�U��   �M�%����]� �����U��Q�M��EP�M��?������؋�]� �U��Q�M��E�3Ƀ8������]���������U��Q�M��E��8�u�M��    �U��E�Z�#�E��8 u�M��A�E������D{	�U��   ��]� ����U��Q�M��E��8�u4�M��    �U����E��M�J�E�B�M�J�E�B�M�J�(�U��: u �EP�M���Q�%   ����t	�U��   ��]� ���������������U��Q�E�M� �������Dz3�U�E�B�@������Dz�M�U�A�B������Dz	�E�    ��E�   �E���]���������U��Q�M��E�����]����������������U��Q�M��E��8�u(�M��    �U����E��M�J�E�B�M�J�(�U��: u �EP�M���Q�!   ����t	�U��   ��]� �����������U����E�M� �������Dz�U�E�B�@������Dz3��T�M�U��J���$�X������E�M� �I���$�]��<������E�������D{	�E�   ��E�    �E��]�������U��Q�M��M��$���E�P�p3�Q$�BD�Ѓ��E���]������U��Q�M��M���#���E�P�p3�Q$�BD�Ѓ��MQ�U�R�p3�H$�Qd�҃��E���]� �����������U��Q�M��M��#���E�P�p3�Q$�BD�Ѓ��MQ�U�R�p3�H$�Q�҃��E���]� �����������U��Q�M��M��A#���E�P�p3�Q$�BD�Ѓ��M�Q�UR�p3�H$�QL�҃��E���]� �����������U��Q�M��E�P�p3�Q$�BH�Ѓ��M��,!����]���������U��Q�M��EP�M�Q�p3�B$�HL�у���]� ����������U��Q�M��EP�MQ�UR�EP�p3�Q$�M��B�Ћ�]� ��U��Q�M��EP�p3�Q$�M��Bl�Ћ�]� ��������������U��Q�M��p3�P$�M��Bp�Ћ�]������U��Q�M��E�P�p3�Q$�B�Ѓ���]�U����M�E�P�M�Q�p3�B$�H�у�P�M��!���M�� ���E��]� ����U��Q�M��EP�M�Q�p3�B$�H�у���]� ����������U��� �M��E�P�M�Q�p3�B$�H �у�P�M�����M��]����E��]� ����U��� �M��E�P�M�Q�p3�B$�H$�у�P�M������M������E��]� ����U��� �M��EP�M�Q�M�������������M�������E��]� ���������������U��Q�M��E�P�p3�Q$�B(�Ѓ���]�U��Q�M��E�P�p3�Q$�Bh�Ѓ���]�U��Q�M��EP�M�Q�p3�B$�H,�у���]� ����������U��Q�M��EP�M�Q�p3�B$�H0�у���]� ����������U����M�E�P�M�Q�p3�B$�Ht�у�P�M�% ���M��M���E��]� ����U��Q�M��EP�M�Q�p3�B$�H4�у���]� ����������U��Q�M��EP�M�Q�p3�B$�H8�у���]� ����������U��Q�M��E�P�MQ�p3�B$�HL�у��E���]� �������U����EP�M�������MQ�U�R�p3�H$�Q@�҃��E�P�M������M��"����E��]������������U��Q�M��EP�M�Q�p3�B$�H@�у��E���]� �������U��Q�M��EP�M�Q�p3�B$�H<�у���]� ����������U��Q�M��EP�M�Q�p3�B$�H<�у��������]� ���U��Q�M��EP�MQ�U�R�p3�H$�QP�҃���]� �������U��Q�M��EP�M�Q�p3�B$�HT�у���]� ����������U��p3�H$�QX��]���������������U��EP�p3�Q$�B\�Ѓ�]�������U��Q�M��EP�MQ�UR�E�P�p3�Q$�B`�Ѓ���]� ��U��p3�H(���]����������������U��E�Q�p3�B(�H�у��U�    ]������������U��Q�M��EP�MQ�UR�EP�MQ�UR�p3�P(�M��B�Ћ�]� �����������U��Q�M��p3�P(�M��B�Ћ�]������U��Q�M��EP�p3�Q(�M��B�Ћ�]� ��������������U��Q�M��EP�MQ�UR�p3�P(�M��B�Ћ�]� �������U��Q�M��EP�MQ�p3�B(�M��P �ҋ�]� ����������U��Q�M�j�EP�MQ�p3�B(�M��P�ҋ�]� ��������U��Q�M��EP�MQ�UR�p3�P(�M��B$�Ћ�]� �������U��Q�M��p3�P(�M��B(�Ћ�]������U��Q�M��p3�P(�M��B,�Ћ�]������U��Q�M��p3�P(�M��B0�Ћ�]������U��Q�M��EP�p3�Q(�M��B4�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M��BX�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M��B\�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M��B`�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M��Bd�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M��Bh�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M��Bl�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M��Bx�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q(�M��Bt�Ћ�]� ��������������U��Q�M��EP�p3�Q(�M��Bp�Ћ�]� ��������������U����M��EP�M�������t/�M��Q�M�������t�U��R�M�������t	�E�   ��E�    �E���]� ��������U����M��EQ� �$�M��F  ��t5�MQ�A�$�M��0  ��t�UQ�B�$�M��  ��t	�E�   ��E�    �E���]� �������������U����M��EP�M�������t/�M��Q�M�������t�U��R�M�������t	�E�   ��E�    �E���]� ��������U����M��E��� �$�M��D  ��t9�M���A�$�M��,  ��t!�U���B�$�M��  ��t	�E�   ��E�    �E���]� �������U����M��EP�M��K�����tB�M��Q�M��8�����t/�U��R�M��%�����t�E��$P�M�������t	�E�   ��E�    �E���]� �����U����M��EP�M��;�����tB�M��Q�M��(�����t/�U��R�M�������t�E��$P�M�������t	�E�   ��E�    �E���]� �����U����M��EP�M��;�����tB�M��Q�M��(�����t/�U��0R�M�������t�E��HP�M�������t	�E�   ��E�    �E���]� �����U����M��EP�M��+�����tB�M��Q�M�������t/�U��0R�M�������t�E��HP�M��������t	�E�   ��E�    �E���]� �����U����M��E�    �E�    �E�P�M��]�����u3��   �}� u#�M����P�M����M��C���   �   h�hj  �M�Q�p3�B���   �у��E��}� uj��M�����3��Lj �U�R�E�P�M��������u�M�Q�1C����3��&j �U���R�E�P�M�  �M�Q�C�����   ��]� ��������������U����M�M��?���E�P�M��������u�E�    �M��p���E���M�Q�M�O����E�   �M��P���E��]� �������U����M��E�P�M��[�����u3���M�����ًU�
�   ��]� ���������U��Q�M��} ����Q�M��  ��]� U����M�j �M��  ���E�h<�h�  �E�P�p3�Q���   �Ѓ��E�}� uj��M�����3��[j �M�Q�U�R�M��  �E�P�M��P  ��t�M�Q�U�R�M��l�����t	�E�   ��E�    �E�E��M�Q�A�����E���]� �������������U����M�E�P�M����P�M��"����E��M������E���]� ��������������U��Q�M��EP�p3�Q(�M��B8�Ћ�]� �������������U��Q�M��EP�p3�Q(�M��B<�Ћ�]� �������������U��Q�M��EP�p3�Q(�M��B@�Ћ�]� �������������U��Q�M��EP�p3�Q(�M��BD�Ћ�]� �������������U��Q�M��EP�p3�Q(�M��BH�Ћ�]� ��������������U��Q�M��EP�MQ�p3�B(�M��P|�ҋ�]� ����������U��Q�M��EP�p3�Q(�M��BL�Ћ�]� ��������������U��Q�M��EP�MQ�p3�B(�M����   �ҋ�]� �������U��Q�M����E�$�p3�P(�M��BT�Ћ�]� ����������U��Q�M�Q�E�$�p3�P(�M��BP�Ћ�]� ������������U��p3�H(�Q��]���������������U��E�Q�p3�B(�H�у��U�    ]������������U��Q�M��E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP�p3�Q(�M����   �Ћ�]�( �������U��EP�MQ�UR�EP�MQ�p3�B(�H�у�]�������U��p3�H,�Q,��]���������������U��Q�M��p3�P,�M��B4�Ћ�]������U��E�Q�p3�B,�H0�у��U�    ]������������U��Q�M��p3�P,�M��B8�Ћ�]������U��� �M��E�P�p3�Q,�M��B<��P�M������M��!����E��]� ��������U����M�EP�M�Q�p3�B,�M�P@��P�M����M��-���E��]� ����U��j j �p3�H,��҃�]���������U��Q�M��EP�MQ�U�R�p3�H,�Q�҃���]� �������U��E�Q�p3�B,�H�у��U�    ]������������U��Q�M��p3�P,�M��B�Ћ�]������U��Q�M��p3�P,�M��B�Ћ�]������U��Q�M��p3�P,�M��B�Ћ�]������U��Q�M��p3�P,�M��B �Ћ�]������U��Q�M��p3�P,�M��B$�Ћ�]������U��Q�M��p3�P,�M��B(�Ћ�]������U��Q�M��EP�MQ�p3�B,�M��P�ҋ�]� ����������U��� �M��E�P�p3�Q,�M��B��P�M������M��1����E��]� ��������U��EP�MQ�UR�p3�H��D  �҃�]�������������U��EP�MQ�UR�p3�H��H  �҃�]�������������U��EP�p3�Q��L  �Ѓ�]����U��EP�MQ�p3�B�H�у�]���U��EP�MQ�UR�p3�H�Q�҃�]����������������U��EP�MQ�p3�B�H�у�]���U��EP�MQ�UR�p3�H�Q�҃�]����������������U��EP�MQ�p3�B�H�у�]���U��EP�MQ�p3�B���  �у�]����������������U��EP�p3�Q�B�Ѓ�]�������U���,�E�P�M������M��V�����u�E�    �M��c����E��~j�M�Q��������u$�U�R��������u�E�    �M��-����E��Hj�EP�}�������u$�MQ�]�������u�E�    �M�������E���E�   �M�������Eԋ�]�������������U��EP�p3�Q�B �Ѓ�]�������U��EP�MQ�p3�B�H(�у�]���U��EP�MQ�UR�EP�MQ�p3�B��  �у�]����U��EP�MQ�UR�EP�p3�Q��   �Ѓ�]��������U��EP�p3�Q��  �Ѓ�]����U��EP�MQ�UR�p3�H��  �҃�]�������������U����E�P�p3�Q�B$�Ѓ�P�M�l����M������E��]��������������U����E�P�p3�Q���  �Ѓ�P�M�)����M��q����E��]�����������U��EP�MQ�p3�B���  �у�]����������������U���D�E�    �=�3 t�E�P��3�{����M��E���M�������M��E��M��M��U�R�M�����E���t�e���M�������M���t�e���M������E��]���U����EP�M�Q�p3�B���  �у�P�M�5����M��}����E��]�������U��j�EP�������E]�����������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��p3�H���   ��]������������U��EP�p3�Q���   �Ѓ��M�    ]�����������U��Q�M��EP�MQ�UR�EP�p3�Q�M���Ћ�]� ���U��Q�M��p3�P�M��B�Ћ�]������U��Q�M��p3�P�M����   �Ћ�]���U��Q�M��EP�p3�Q�M��B`�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��Bd�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��Bh�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��Bl�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��Bp�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��Bt�Ћ�]� ��������������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M���  �Ћ�]� �����������U��Q�M��EP�p3�Q�M��Bx�Ћ�]� ��������������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M��B|�Ћ�]� ��������������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�M�Q�p3�B��  �у���]� �������U��Q�M��EP�MQ�p3�B�M����   �ҋ�]� �������U��Q�M��EP�MQ�p3�B�M����   �ҋ�]� �������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U����M��} t&�EP�M�Q�p3�B �H$�у���t	�E�   ��E�    �E���]� �����������U��Q�M��E�P�MQ�UR�p3�H �QL�҃���]� �������U��Q�M��} u3���EP�M�Q�p3�B �H(�у��   ��]� �����������U��Q�M��EP�p3�Q�M��B�Ћ�]� �������������U��Q�M��EP�p3�Q�M��B�Ћ�]� �������������U��Q�M��EP�p3�Q�M��B�Ћ�]� �������������U��Q�M��EP�p3�Q�M��B�Ћ�]� �������������U��Q�M��EP�p3�Q�M��B�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��B�Ћ�]� ��������������U��Q�M��EP�MQ�p3�B�M��P\�ҋ�]� ����������U��Q�M��EP�MQ�p3�B�M���  �ҋ�]� �������U��Q�M����E�$�p3�P�M��B �Ћ�]� ����������U��Q�M�Q�E�$�p3�P�M��B$�Ћ�]� ������������U��Q�M����E�$�p3�P�M��B(�Ћ�]� ����������U��Q�M��EP�p3�Q�M��B,�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��B0�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��B4�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��B8�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��B<�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��B@�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��BD�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��BH�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��BL�Ћ�]� ��������������U��Q�M��EP�p3�Q�M��BP�Ћ�]� ��������������U��Q�M��EP�MQ�UR�EP�p3�Q�M����   �Ћ�]� ���������������U��Q�M��EP�p3�Q�M��BT�Ћ�]� ��������������U��Q�M��EP�M�Q�p3�B��  �у���]� �������U��Q�M��EP�MQ�UR�EP�p3�Q�M����   �Ћ�]� ���������������U��Q�M��EP�MQ�UR�EP�p3�Q�M����   �Ћ�]� ���������������U��Q�M��EP�MQ�p3�B�M��PX�ҋ�]� ����������U��Q�M��p3�P�M����   �Ћ�]���U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U��Q�M��EP�MQ�p3�B�M����   �ҋ�]� �������U��Q�M��p3�P�M����   �Ћ�]���U��Q�M��EP�MQ�p3�B�M����   �ҋ�]� �������U��Q�M��p3�P�M����   �Ћ�]���U��Q�M��p3�P�M����   �Ћ�]���U��Q�M��p3�P�M����   �Ћ�]���U��EP�MQ�UR�EP�MQ�p3�B���   �у�]����U��EP�MQ�UR�EP�p3�Q��   �Ѓ�]��������U����EP�MQ�U�R�p3�H���  �҃�P�M�"����M��J����E��]����U��EP�MQ�p3�B���  �у�]����������������U��Q�M��EP�MQ�UR�E�P�p3�Q�B�Ѓ���]� ��U��Q�M��EP�p3�Q�M��Bd�Ћ�]� ��������������U��Q�M��EP�MQ�UR�p3�P�M��Bh�Ћ�]� �������U��� �M�j h�  �M��X  �} u�   �kj h�  �M���  �E��}� u3��O�M���P  �EPh�  �M��������E�$h�  �M������j �M�Q�M��-  �E�   �M��CQ  �E��]� ����������U��Q�M����E�$�E�P�p3�QH�B�Ѓ���]� �����U��Q�M��EP�M�Q�p3�BH���   �у���]� �������U��Q�M��EP�M�Q�p3�BH���  �у���]� �������U��Q�M��EP�M�Q�p3�BH���  �у���]� �������U��Q�M��EP�MQ�U�R�p3�HH��  �҃���]� ����U��Q�M��EP�MQ�U�R�p3�HH��  �҃���]� ����U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��Q�M��EP�M�Q�p3�BH���  �у���]� �������U��Q�M�j �E�P�p3�QH���   �Ѓ���]������������U��Q�M��EPj �M�Q�p3�BH���   �у���]� �����U��Q�M�j�E�P�p3�QH���   �Ѓ���]������������U��Q�M��EPj�M�Q�p3�BH���   �у���]� �����U��Q�M�j�E�P�p3�QH���   �Ѓ�����؋�]������U��Q�M��EPj�M�Q�p3�BH���   �у���]� �����U��Q�M��EP�MQ�U�R�p3�HH���   �҃���]� ����U��Q�M��EP�MQ�U�R�p3�HH���   �҃���]� ����U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�HH���  �҃���]� ��������U����M��EP��  ���E��}� t�MQ�U�R�M������E���]� ���������U����M��EP�MQ�*�  ���E��}� t�UR�E�P�M������E���]� �����U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��Q�M��EP�M�Q�p3�BH���   �у���]� �������U��Q�M��EP�MQ�U�R�p3�HH���  �҃���]� ����U��Q�M��EP�M�Q�p3�BH���   �у���]� �������U��Q�M��EP�MQ�U�R�p3�HH��8  �҃���]� ����U��Q�M��EP�MQ�U�R�p3�HH��   �҃���]� ����U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��Q�M��E�P�p3�QH��  �Ѓ���]��������������U��Q�M��E�P�p3�QH��  �Ѓ���]��������������U��Q�M��EP�MQ�U�R�p3�HH��  �҃���]� ����U��Q�M��EP�MQ�UR�E�P�p3�QH��   �Ѓ���]� ���������������U��Q�M��EP�MQ�UR�EP�M�Q�p3�BH��|  �у���]� �����������U��Q�M��EP�M�Q�p3�BH��  �у���]� �������U��Q�M��E�P�p3�QH��T  �Ѓ���]��������������U��Q�M��EP�MQ�U�R�p3�HH��  �҃���]� ����U��Q�M��EP�M�Q�p3�BH��8  �у���]� �������U��Q�M��EP�M�Q�p3�BH��<  �у���]� �������U��Q�M��EP�MQ�UR�E�P�p3�QH��@  �Ѓ���]� ���������������U��Q�M��EP�M�Q�p3�BH���  �у���]� �������U��Q�M��E�P�p3�QH��L  �Ѓ���]��������������U��Q�M��EP�M�Q�p3�BH��H  �у���]� �������U����M�j h�  �M���$  �������E��M���$  ���}�u�E���3���]���������������U��Q�M�j h�  �M���������������]����������������U����M�EP�MQ���E�$�U�R�E�P�p3�QH��  �Ѓ��M���P�Q�P�Q�P�Q�P�Q�@�A�E��]� ������������U����M�EP�MQ���E�$�U�R�E�P�p3�QH��  �Ѓ��M���P�Q�P�Q�P�Q�P�Q�@�A�E��]� ������������U��Q�M��EP�MQ�UR�E�P�p3�QH��   �Ѓ���]� ���������������U��p3�HH��  ��]������������U��EP�p3�QH��  �Ѓ�]����U��Q�M����E�$�E�P�p3�QH��$  �Ѓ���]� ��U��Q�M��E�P�p3�QH��(  �Ѓ���]��������������U��Q�M��EP�MQ�U�R�p3�HH��,  �҃���]� ����U��Q�M��EP���E�$�MQ�U�R�p3�HH��0  �҃���]� �����������U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��Q�M��E�P�p3�QH��4  �Ѓ���]��������������U��Q�M��E��     �E���]����������U��Q�M�j�E��Q�p3�BH��|  �у���]����������U��Q�M��EP�p3�QH��x  �Ѓ��M���U�3��: ����]� �����������U��Q�M�j �E��Q�p3�BH��|  �у���]����������U��Q�M��E�P�p3�QH��P  �Ѓ���]��������������U��Q�M��E�P�p3�QH��T  �Ѓ���]��������������U��Q�M��E�P�p3�QH��X  �Ѓ���]��������������U����M�E�P�M�Q�p3�BH��\  �у��U��
�H�J�H�J�H�J�H�J�@�B�E��]� �������������U��Q�M��E�P�p3�QH��`  �Ѓ���]��������������U��Q�M��EP�M�Q�p3�BH��d  �у���]� �������U��Q�M����E�$�E�P�p3�QH��h  �Ѓ���]� ��U��Q�M����E�$�E�P�p3�QH��t  �Ѓ���]� ��U��Q�M����E�$�E�P�p3�QH��l  �Ѓ���]� ��U��Q�M��EP�M�Q�p3�BH��p  �у���]� �������U��Q�M��EP�MQ�UR�EP�M�Q�p3�BH���  �у���]� �����������U��Q�M��EP�MQ�UR�EP�MQ�UR�E�P�p3�QH���  �Ѓ���]� ���U��E P�MQ���E�$�UR�EP�MQ�p3�BH���   �у�]�����������U��EP���E�$�MQ�UR�EP�p3�QH���   �Ѓ�]���������������U���E�M�P��L�  �E�EP�MQ�UR�h  ��]����U���   V�M��  �E��E�    �M�  �E��E�    �E�    �E�    �E�    �}� u
�   �E  �M�5  =�  ��  j h:  �M�;  �EЋM�  �E��E�    �M��  �E��M�3  �E��M�  �E��E�    �	�E����E��M�;M���   �}� taj��U�R�M��Ӵ  �E��}��tJ�M�k�M��<  9E�t빋M�k�M����  �E��E�;E�~�M��MȋM�k�M��X�  E�E��0�U����E����M��u��T;Tu�E���E��	�M���M��O����}� tj �UR�M��G�  ��u
��
  ��
  �}� tj�M��k�  ��t^�M��o�  ;E�uQh��h�  �E�k�P�p3�Q���  �Ѓ��E��}� u
�
  �
  �M�Q�U�R�M���  P�!  ��h��h�  �E�k�P�p3�Q���  �Ѓ��E��}� u
�H
  �C
  �M�Q�U�R�E�P��   ���}� ~;h��h�  �M�����Q�p3�B���   �у��E�}� u
��	  ��	  j��U�R�M�������u
��	  ��	  �}� tj�EP�M���  ��u
�	  �	  �}� t�M��P�  ��|����
ǅ|���    ��|����M�M��  �E��E�    �E�    �	�U����U��E�;E���  �}� �4  j��M�Q�M��}�  �E��}���  �M�k�M���  9E�t뱋M�k�M���  �E��E�    �E�    �E�    �	�Uă��UċM�k�M��,���9E��  �E�P�M�k�M��A  ��u�ȋM�Q�M�k�M���  �E��U����EԋM�u�����Eԃ��EԋM����UԋE���Mԃ��MԋU����EԋM�u��T���Eԃ��EԋM���   �EԋM���Uԃ��UԋE����MԋU�u��D���Mԃ��MԋU���   �MԋU���Eԃ��EԋM����UԋE�u��L���Uԃ��UԋE���   �UԋE���Mԃ��M�������UԉU��}� ��  �E��+���P�E�P�M��U  �E�    �M�;M�|
�  �~  �UԋE���M��}� t4�U�k�U��E�k�E�
��J�H�J�H�J�H�J�H�R�P�E�k�E��M�k�M����P�Q�P�Q�P�Q�P�Q�@�A�M�;M���   �UԋE��;M���   �UԋE�D��������E��MԋU�D����E��M���x�����x���wR��x����$��4�E����M��U��4�E����M��U�T�"�E����M��U�T��E����M��U�T�Eԃ��E��J����M���M�U����U��E�;E�������M�;M�t
�#  �  �  �U����E����M��u��T3�;T���M܃}� �  �U����E��k�M��U�k�U���A�B�A�B�A�B�A�B�I�J�U����E��Lk�M��U��k�U���A�B�A�B�A�B�A�B�I�J�U����E��Lk�M��U��k�U���A�B�A�B�A�B�A�B�I�J�}� tA�U����E��Lk�M��U��k�U���A�B�A�B�A�B�A�B�I�J�U����E��k�M��U�k�U����A�B�A�B�A�B�A�B�I�J�U����E��M��U���U�E����M��Tk�U��E�k�E��
��J�H�J�H�J�H�J�H�R�P�E����M��U�T�E���E�M����U��D
k�E��M�k�M����P�Q�P�Q�P�Q�P�Q�@�A�M����U��E�D
�M���M�}� tY�U����E��Lk�M��U�k�U����A�B�A�B�A�B�A�B�I�J�U����E��M�L�U���U���E����M����U��u��D�D
������M�Q�k�����U�R�_�����6  �M�_  =  �#  �M��  �E��M�  �E��E�    �	�E����E��M�;M�}D�U��E��<� u��M��U��|� t�E��M����E�P�M���U��E��ЋU�DJ��E��h �hY  �M�k�Q�p3�B���  �у��E��}� u3��  �U�R�E�P�M�Q�  ��h(�h^  �U���R�p3�H���  �҃��E��}� u3��k  �E�P�M�Q�U�R�"  ���E�+���P�E�P�M�
�����u�M�Q������U�R�����3��  �M�_  �E��M�  �E��E�    �E�    �E�    �	�E����E��M�;M��\  �U��E��<� u���E�    �	�M����M��U����E��M�;���   �U�U�k�U��E�k�E��
��J�H�J�H�J�H�J�H�R�P�E����E��M��U��D
k�E��M�k�M����P�Q�P�Q�P�Q�P�Q�@�A�M����M��Y����U��E��|� t}�M�M�k�M��U�k�U����A�B�A�B�A�B�A�B�I�J�U����U��E�k�E��M�k�M����P�Q�P�Q�P�Q�P�Q�@�A�M����M��U��E��M�ЉM������E�    �	�U����U��E�+���9E�}�E��M��D�    �U��E���   �͍M�Q�$�����U�R������   �&�E�P������M�Q��
�����U�R��
����3�^��]ÍI !.2.D.V.U����M��E�    �E�    �E�    �E�8 u'�MQ�M��~  ��uj�M��@  ��u	�E�    ��E�   �U�E��M�9 uc�M��  �} u�UR�EP�MQ�UR�EP�M��"  �7�M�M���M��  �E�}� t�UR�EP�MQ�U�R�EP�M���  �ыM�9 u�M��I  ��t	�E�    ��E�   �U�E��M�9 u�M��M  �UR�M��A  �   �M���   �} u�EPj �MQ�UR�EP�M��t  �E��uh  �%	  ���E��}� u3��^�M�}  P�M��  �M�M���M��  �E�}� t1�URj �EP�M�Q�UR�M��  �E��}� t�E�P�M���  뾋E���]� �U��Q�M��E�P�MQ�UR�p3�HH���   �҃���]� ����U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��Q�M��EP�MQ�U�R�p3�HH���   �҃���]� ����U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�HH���  �҃���]� ��������U��Q�M��E�P�p3�QH��t  �Ѓ���]��������������U��Q�M��E�� \��M��A    �E���]����������������U��Q�M��E�� \��M��QR�p3�Hl�Q�҃���]������U��Q�M��E��HQ�p3�Bl�H�у��} u�   �1�UR�EP�MQ�UR�p3�Hl��҃��M��A�U�3��z ����]� �������������U��Q�M��E��x u3���M��QR�p3�Hl�Q�҃���]��U����M�E�P�M�Q�UR�EP�M���  �M�;Mu�E����U�;Uu�E�������]� ����������U��EP���E�$�MQ�UR�p3�HH���  �҃�]����U��EP�MQ�UR�EP�p3�QH���  �Ѓ�]��������U��E P�MQ�UR�EP�MQ�UR�EP�p3�QH���  �Ѓ�]������������U��E0P���E(�$�M$Q�U R�EP�MQ�UR�EP�MQ�UR�p3�HH���  �҃�,]������������U��EP�MQ�UR�p3�HH���  �҃�]�������������U��Q�M��EP���E�$�M�Q�p3�BH���  �у���]� ��������������U����M��E�    �}u�M��"����E��$�} u�M�������E���}u�M��,����E��}� u3���E�P�MQ�M��   ��]� ���������U���$V�M�葶  �E�}� t�} u3���   �M���  �E��M��h  ���E��}� u�E���   �E�    �	�E����E��M誶  9E���   �M�Q�U�R�E�P�M�Q�M蹷  ��u�ȋU�U��	�E����E��M�;M�_�U�����u$�E������M������U��u��D;Du���M���Q�M�|  �U����D��E�}��t�M�Q�M��-�  ��K����E�^��]� ������������U���V�M�M���  �E�}� u3��G  �E�    �}u�M��y����E��$�} u�M��6����E���}u�M������E��}� u3���   �M��+�  �E�    �	�E����E��M���
  9E���   �M�Q�M�  �E��}� u�ϋU��BP�M�  ��t�M���Q�M��?�  �U��BP�M�  ��t�M���   R�M���  �E����M����U�u�D;Dt&�M��QR�M�N  ��t�E���   Q�M��״  �U��BP�M�(  ��t�M���   R�M�豴  �����   ^��]� U��E P�MQ�UR�EP�MQ�UR�EP�p3�QH���   �Ѓ�]������������U��Q�M��E�P�p3�QH���   �Ѓ���]��������������U��EP�MQ�UR�EP�MQ�p3�BH���  �у�]����U����E�$���E�$�����$�EP�M�������$�\  ���$�MQ�M�z���]���������U���H�M��2���P�EP�M�Q�M�������E�$���E�$���E��$�  ���$���E�$���E�$���E��$��  ���$���E�$���E�$���E��$�  ���$�M�����P�UR�M�������]�������U��EP�p3�QH��Ѓ�]��������U��E�Q�p3�B@�H�у��U�    ]������������U��h�  �p3�HH��҃�]��������U��E�Q�p3�B@�H�у��U�    ]������������U��Qh  �R������E��}� u3��jj �EPh�  �M�������u�.�,j �MQh(  �M��������u��j j�M���
  �E��#�}� t�U�R�p3�H@�Q�҃��E�    3���]�����U��E�Q�p3�B@�H�у��U�    ]������������U��Qh�  �������E��}� u3��8�EP�MQ�M��������u!�}� t�U�R�p3�H@�Q�҃��E�    �E���]�������U��E�Q�p3�B@�H�у��U�    ]������������U��EP�MQ�p3�BH�H�у�]���U��E�Q�p3�B@�H�у��U�    ]������������U��Q�M��EP�M�Q�p3�BH���  �у���]� �������U��Q�M��EP�M�Q�p3�BH���  �у���]� �������U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��EP�MQ�p3�BH���  �у�]����������������U��E0P�M,Q�U(R�E$P�M Q���E�$���E�$�UR�EP�p3�QH��P  �Ѓ�,]����������U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��Q�M��EP�MQ�U�R�p3�HH���  �҃���]� ����U��Q�M��E�P�p3�QH��  �Ѓ���]��������������U��Q�M��EP�MQ�UR�E�P�p3�QH���  �Ѓ���]� ���������������U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��Q�M��E�P�p3�QH���  �Ѓ���]��������������U��Q�M��EP�M�Q�p3�BH��  �у���]� �������U��Q�M��EP�M�Q�p3�BH��  �у���]� �������U��Q�M��E���]���U��Q�M���]������U��p3�HH���  ��]������������U��EP�p3�QH���  �Ѓ�]����U��Q�M��E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R�p3�HH���  �҃�0��]�, U��Q�M��E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R�p3�HH���  �҃�0��]�, U��Q�M��E�P�p3�QH��,  �Ѓ���]��������������U��Q�M��EP�M�Q�p3�BH��X  �у���]� �������U��Q�M��E�P�p3�QH��\  �Ѓ���]��������������U��EP�MQ�UR�EP�MQ�p3�BH��0  �у�]����U��Q�M��EP�MQ�U�R�p3�H@�Q(�҃���]� �������U��Q�M��E�P�p3�Q@�B,�Ѓ���]�U��Q�M�h�  �M��   ��]���������U��Q�M��EP�M�Q�p3�BH���   �у���]� �������U��E;E}�E��M;M~�E��E]���������������U��Q�M��p3���   �M��B�Ћ�]���U��Q�M��EP�MQ�U�R�p3�HH���   �҃���]� ����U��Q�M�j h�  �M��
   ��]�������U��Q�M��EP�MQ�U�R�p3�HH���   �҃���]� ����U��Q�M�j h(  �M�������]�������U��Q�M�h(  �M��������]���������U��Q�M�j h�  �M��z�����]�������U��Q�M�h�  �M�������]���������U��Q�M��E���U���	   ��]� ���U��Q�M��E�� %�������]���������U��Q�M��E���U���	   ��]� ���U��Q�M��E�� %   ��������]�����U����M��E��x ~�M��	�����E���E������E���]��U��Q�M��EP�p3���   �M��BH�Ћ�]� �����������U��Q�M��p3���   �M��Bx�Ћ�]���U��Q�M��EP�p3���   �M��B|�Ћ�]� �����������U��Q�M��p3���   �M��B(�Ћ�]���U��Q�M��EP�M�Q�p3�BH���   �у���]� �������U��Q�M��EP�M�Q�p3�BH���   �у���]� �������U��Q�M��EP�M�Q�p3�BH���   �у���]� �������U��Q�M��M��a����E��t�M�Q��������E���]� ����U��Q�M��EP�MQ�UR�EP�M��QR�p3�Hl�Q�҃���]� ������������U��Q�M�j h�  �M��
   ��]�������U��Q�M��EP�MQ�U�R�p3�HH��p  �҃���]� ����U��Q�M��EP�M��QR�p3�Hl�Q�҃���]� ��������U��Q�M��EP�M�Q�p3�B\�H,�у���]� ����������U���E�]����Au�E��E�]����z�E��E]�����U��Q�M��EP�MQ�p3���   �M��P�ҋ�]� �������U��Ek�P�MQ�UR詹  ��]�����U��Q�M��}~�EP�MQ�UR�M��/   ��]� ���������U��E��P�MQ�UR�Y�  ��]�����U����M�E�M���U��EP�M��?   ��P�M�Q�UR�E�P�M��h   �MQ�U�R�EP�M�Q�M��  ��]� ����������U����M��E�    ��E���E�}t�M����M���E���]� ������������U����M�E+E���� ��   �} u�MQ�UR�EP�M��  �v�M���M�U��R�E+E���+����M��R�EP�MQ�M���   �E��U�R�EP�MQ�UR�M��Y  �E��EP�MQ�U�R�EP�M��^����M��M�\�����]� �������������U����M��} ~5�E   �E��M�Q�UR�EP�M��  �MQ�U�R�EP�M��  ��M;Mt�UR�EP�MQ�M���   ��]� ����������U��Q�M��EP�MQ�   ����t;�UR�EP�x   ����t�E�Y��MQ�UR�]   ����t�E�>�E�9�4�EP�MQ�=   ����t�E���UR�EP�"   ����t�E��E��]� �������������U��E�M�3�;��]�������������U����p!3ŉE��M�E+E���� ~�M+M��Q�UR�EP�M���  �   �M���M��U��U�E���E���M���M�U����U��E�;EtL�M�Q�U�R�_�������t8j�E�P�M�Q�)�  ��j�U�R�E�P��  ��j�M�Q�U�R��  ��뚋E����E��M�;M�t����M�3��B�  ��]� �����������U����p!3ŉE��M��E���E�   ����   �U���U�EP�MQ��������t��U���U�EP�MQ��������t��U;Ur�E�Yj�EP�M�Q�M�  ��j�UR�EP�;�  ��j�M�Q�UR�)�  ���E;Eu�M�M��U;Uu�E�E�O����M�3��Z�  ��]� ���U��Q�M��	�E���E�M;Mt�UR�EP�M��  �݋�]� ��������������U���,�p!3ŉE�Mԃ}}�Z  �E�E��E��+������E��   ���9  �}�~�U����U��c�E����E��M��U�D���E܋M��U�ʉE�j�M�Q�U�R�/�  ��j�E�P�M�Q��  ��j�U�R�E�P��  ���}���   �M��M�U�E�L���M�U���;U���   �E�E؋M���M�U�E�L���M�U�;U�})�E��P�M�Q���������t�U���U�E���E�M�Q�U�R��������t8j�E�P�M�Q�m�  ��j�U�R�E�P�[�  ��j�M�Q�U�R�I�  �����S��������M�3�菶  ��]� ��������U����p!3ŉE��M�E��P�MQ��������t_j�UR�E�P��  ���M��M�j�U��R�EP�̲  ���M���M�U��R�E�P���������u�j�M�Q�UR蚲  ���M�3���  ��]� �������U����M��E�M��;t3���   �E�x uE�M�9 u=�U�z u4�E��x u�M��9 u�U��z u	�E�   ��E�    �E��   �I�E��x u@�M��9 u8�U��z u/�E�x u�M�9 u�U�z u	�E�   ��E�    �E��M�E�x t�M��y t�U�E��J;Ht3��)�U�z t�E��x t�M�U��A;Bt3���   ��]� ����������U��Q�M��EP�M�������������]� U����M��E�    �	�E����E��M�Q�M���  �8 t��E���]������������U����M��E�    �	�E����E��M�Q�M��  �8 t(�U�R�M�x  P�E�P�M��k  ���T�����t�뾃} t�M�U���}� ~�E�P�M��<  �8 u	�E�   ��E�    �E��]� ��������������U��Qj�5   ���E��}� t	�E��x u3���MQ�UR�EP�M��Q�҃���]��U��hx3�EPhD �Z�  ��]������U����M�j\��������E��}� t	�E��x\ u��M�Q�U��B\�Ѓ��E���]����U����M�j\�������E��}� t	�E��x\ u��M�Q�U��B\�Ѓ��MQ�M���  �E���]� �����U����M�j\�@������E��}� t	�E��x\ u��M�Q�U��B\�Ѓ��MQ�M��~  �E���]� �����U����M�j\��������E��}� t	�E��x\ u�$�M�Q�U��B\�Ѓ��MQ�M��  P�M��%  �E��]� ������������U����M�j\�������E��}� t	�E��x\ u�'�M�Q�U��B\�Ѓ��MQ�M���   �UR�M��  �E���]� ���������U����M�j\�0������E��}� t	�E��x\ u�3�M�Q�U��B\�Ѓ��MQ�M��n   �UR�M��   �EP�M��   �E���]� �������������U����M�j`��������E��}� t	�E��x` u��M�Q�U��B`�Ѓ���]�������U����M�jd�������E��}� t	�E��xd u��MQ�U�R�E��Hd�у���]� U����M�jh�@������E��}� t	�E��xh u��MQ�U�R�E��Hh�у���]� U����M�jl� ������E��}� t	�E��xl u��M�Q�U��Bl�Ѓ���]�������U����M�h�   �������E��}� t�E����    u3���MQ�U�R�E����   �у���]� �����U����M�h�   �m������E��}� t�E����    u3���MQ�U�R�E����   �у���]� �����U����M�jp� ������E��}� t	�E��xp u�|3��MQ�U�R�E��Hp�у���]� �����������U����M�jt��������E��}� t	�E��xt uh|3�M�^����E�+�MQ�U�R�E�P�M��Qt�҃�P�M������M������E��]� ��������U����M�jx�`������E��}� t	�E��xx u�E���M�Q�UR�E��Hx�у��E���]� ����������U����M�j|�������E��}� t	�E��x| u3���M�Q�UR�E��H|�у���]� ��������������U����M�j|��������E��}� t	�E��x| u�   ��M�Q�UR�E��H|�у��������]� ����U����M�h�   �m������E��}� t�E����    u�E��%�MQ�U�R�E�P�M����   �҃��M��^����E���]� �����U��Q�M��E���]���U��Qj�������E��}� t	�E��x u3���M��Q�ҋ�]�U��Q�E�8 u�6j��������E��}� t	�M��y u��UR�E��H�у��U�    ��]���������U����M��} u3��7j�v������E��}� t	�E��x u3���MQ�UR�E�P�M��Q�҃���]� U����M�j�0������E��}� t	�E��x u3���MQ�U�R�E��H�у���]� ��������������U����M�j��������E��}� t	�E��x u3���MQ�U�R�E��H�у���]� ��������������U����M�j �������E��}� t	�E��x  u3���M�Q�U��B �Ѓ���]�����U����M�j$�P������E��}� t	�E��x$ u3���M�Q�U��B$�Ѓ���]�����U����M�j(�������E��}� t	�E��x( u3���MQ�UR�EP�M�Q�U��B(�Ѓ���]� ������U����M�j,��������E��}� t	�E��x, u3���MQ�UR�E�P�M��Q,�҃���]� ����������U����M�j(�p������E��}� t	�E��x0 u3���MQ�UR�EP�M�Q�U��B0�Ѓ���]� ������U����M�j4� ������E��}� t	�E��x4 u3���M�Q�U��B4�Ѓ���]�����U����M�j8��������E��}� t	�E��x8 u3���MQ�UR�EP�MQ�U�R�E��H8�у���]� ��U����M�j<�������E��}� t	�E��x< u��MQ�U�R�E��H<�у���]� U����M�jD�P������E��}� t	�E��xD u3���M�Q�U��BD�Ѓ���]�����U����M�jH�������E��}� u��EP�M�Q�U��BH�Ѓ���]� ���������U����M�jL��������E��}� u3���EP�M�Q�U��BL�Ѓ���]� �������U����M�jP�������E��}� u3���EP�MQ�U�R�E��HP�у���]� ���U����M�jT�P������E��}� u3���E�P�M��QT�҃���]��������������U����M�jX�������E��}� u��EP�M�Q�U��BX�Ѓ���]� ���������U����M�h�   ��������E��}� u3��&�EP�MQ�UR�EP�MQ�U�R�E����   �у���]� �U����M�h�   �}������E��}� u3���EP�MQ�UR�E�P�M����   �҃���]� ���������U����M�h�   �-������E��}� u3���EP�M�Q�U����   �Ѓ���]� �U����M�h�   ��������E��}� u3���EP�M�Q�U����   �Ѓ���]� �U����M�h�   �������E��}� u3���EP�M�Q�U����   �Ѓ���]� �U����M�h�   �m������E��}� u��EP�MQ�UR�E�P�M����   �҃���]� �����������U���h�   � ������E��}� u�M�L����E�*�EP�M�Q�U����   �Ѓ�P�M�H����M��p����E��]����������U���h�   ��������E��}� t�E����    u�MQ�M������E�.�UR�EP�M�Q�U����   �Ѓ�P�M������M������E��]������U����M�h�   �M������E��}� t�E����    uj �M��  P�M������E�*�MQ�U�R�E��M䋐�   ��P�M�^����M��&����E��]� �������������U����M�h�   ��������E��}� t�E����    u3���MQ�UR�EP�U��M����   �Ћ�]� �U����M�h�   �}������E��}� t�E����    u3���MQ�U��M����   �Ћ�]� ���������U����M�h�   �-������E��}� t�E����    u3���MQ�U��M����   �Ћ�]� ���������U����M�h�   ��������E��}� t�E����    u3���MQ�U��M����   �Ћ�]� ���������U����M�h�   �������E��}� t�E����    u3���U��M����   �Ћ�]����������������U����M�h�   �=������E��}� t�E����    u3���MQ�UR�EP�U��M����   �Ћ�]� �U����M�h�   ��������E��}� t�E����    u��MQ�U��M����   �Ћ�]� �����������U����M�h�   �������E��}� t�E����    u3���MQ�UR�EP�U��M����   �Ћ�]� �U����M�h�   �M������E��}� t�E����    u3���U��M��   �ЉE��E���]����������U��Q�M��E��M��U��B    �E��@    �E���]� ����U��Qj�E   ���E��}� t	�E��x u����'�M Q�UR�EP�MQ�UR�EP�MQ�U��B�Ѓ���]�U��h�3�EPh�f ��  ��]������U���j��������E��}� t	�E��x u�E������M�����E��?�M8Q�U4R�E0P�M,Q�U(R���̍EP�����MQ�U��B�Ѓ�4�E�M�>����E��]��������U��Qj�U������E��}� t	�E��x u3���MQ�UR�E��H�у���]������U��Qj�������E��}� t	�E��x u3���MQ�U��B�Ѓ���]����������U����M��E�P�p3���   �BX�Ѓ��E��}� u3���MQ�UR�M��"  ��]� ������������U����M��E�P�p3���   �BX�Ѓ��E��}� u3���MQ�UR�M��  ��]� ������������U��Q�M��E��M�j j j �U��P�p3�Q�B�Ѓ��M��A�E���]� �����U��Q�M�j j j �E��Q�p3�B�H�у��U��B��]���U��Q�M��E��x u3��1�M��QR�EP�MQ�U��P�p3�Q�B�Ѓ��M��A�   ��]� �����U��Q�M��EP�MQ�U�R�p3�H|�Q�҃���]� �������U��Q�M��EP�MQ�U�R�p3�H|�Q8�҃���]� �������U��Q�M�j j��p3�P�M��B�ЋE���]���������������U��Q�M�j �EP�p3�Q�M��B�ЋE���]� ���������U��Q�M��EPj��p3�Q�M��B�ЋE���]� ���������U��Q�M��M���  ��]��������������U��Q�M�j j �E�P�M�  �E���]� U��Q�M��EP�M�Q�p3�B�H�у���]� ����������U��Q�M��EP�M�Q�p3�B�H�у��������]� ���U����M��EP�M��  �E��M��`  ��]� ����������U��Q�M�h#  �EP�MQ�M��  ��]� ��������������U��Q�M�hF  �EP�MQ�M��d  ��]� ��������������U����M��EP�M��  �E��MQ�M��\  ��]� ������U��Q�M��EP�p3�Q�M����   �Ћ�]� �����������U����M��EP�p3�Q�M����   �ЉE��}� u3���M��
{����]� ����U��Q�M��p3�P�M��B�Ћ�]������U��Q�M��EP�MQ�UR�p3�P�M����   �Ћ�]� ����U��Q�M��E�P�p3���   �BX�Ѓ���]��������������U��Q�M��EP�p3�Q�M��Bt�Ћ�]� ��������������U��Q�M��EP�MQ�UR�p3�P�M��Bl�Ћ�]� �������U��Q�M��EP�M�Q�p3���   �H`�у���]� �������U��Q�M��EP�M�Q�p3�B8�HD�у���]� ����������U��p3�H8�Q<��]���������������U��E�Q�p3�B8�H@�у��U�    ]������������U��p3�H8���]����������������U��E�Q�p3�B8�H�у��U�    ]������������U��Q�M��EP�MQ�UR�E�P�p3�Q8�B�Ѓ���]� ��U��Q�M��EP�MQ�U�R�p3�H8�Q�҃���]� �������U��Q�M��E�P�p3�Q8�B�Ѓ���]�U��Q�M��EP�M�Q�p3�B8�H �у���]� ����������U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�H8�Q$�҃���]� �����������U��Q�M��EP�MQ�UR�EP�MQ�UR�E�P�p3�Q8�B�Ѓ���]� ������U��Q�M��EP�MQ�U�R�p3�H8�Q(�҃���]� �������U��Q�M��EP�MQ�UR�E�P�p3�Q8�B,�Ѓ���]� ��U��Q�M��EP�MQ�UR�E�P�p3�Q8�B�Ѓ���]� ��U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�H8�Q�҃���]� �����������U��Q�M��EP�MQ�U�R�p3�H8�Q0�҃���]� �������U��Q�M��EP�MQ�UR�E�P�p3�Q8�B4�Ѓ���]� ��U��Q�M��EP�M�Q�p3�B8�H8�у���]� ����������U��EP�MQ�UR�EP�p3�Q��x  �Ѓ�]��������U��EP�MQ�p3�B��|  �у�]����������������U��EP�MQ�p3�B���  �у�]����������������U��EP�MQ�p3�B���  �у�]����������������U��EP�p3�Q���  �Ѓ�]����U��EP�p3�Q�B,�Ѓ�]�������U��E P�MQ�UR�EP�MQ�UR�EP�p3�Q���  �Ѓ�]������������U����M��Ҡ���E�P�p3�Q�B8�Ѓ��M�Q�M�Ѡ���M�������E��]���U��p3�H�Q<��]���������������U��EP�MQ�p3�B�H@�у�]���U��p3�H�QD��]���������������U��p3�H�QH��]���������������U��EP�MQ�UR�p3�H�QL�҃�]����������������U��EP�MQ�p3�B�HP�у�]���U��EP�p3�Q��<  �Ѓ�]����U��EP�p3�Q��,  �Ѓ�]����U��E��PP�M��@Q�U��0R�E�� P�M��Q�UR�EP�p3�Q���   �Ѓ�]�������������U��p3�H���   ��]������������U��p3�H���  ��]������������U��EP�MQ�UR�EP�MQh�6  �p3�B���   �у�]���������������U��EP�p3�Q�B�Ѓ�]�������U��EP�p3�Q��\  �Ѓ�]����U��� �EPj hd��M��w���P�M�Q��u�����M�袜���U�R�p3�H�Q�҃��M�膜����]���U��EP�p3�Q�BT�Ѓ�]�������U��EP�p3�Q�BX�Ѓ�]�������U��EP�p3�Q�B\�Ѓ�]�������U��p3�H�Q`��]���������������U��EP�p3�Q���  �Ѓ�]����U��p3�H�Qd��]���������������U��p3�H�Qh��]���������������U��EP�p3�Q�Bl�Ѓ�]�������U��EP�p3�Q�Bp�Ѓ�]�������U��EP�MQ�UR�p3�H�Qt�҃�]����������������U��EP�p3�Q��D  �Ѓ�]����U��EP�MQ�UR�EP�p3�Q��  �Ѓ�]��������U��EP�MQ�p3�B�Hx�у�]���U��EP�MQ�p3�B��@  �у�]����������������U����M��x���E�P�MQ�p3�B�H|�у��U�R�M�x���M��y���E��]���������������U��EP�MQ�p3�B���   �у�]����������������U��EP�MQ�p3�B��h  �у�]����������������U��EP�MQ�UR�EP�p3�Q��d  �Ѓ�]��������U��EP�MQ�UR�p3�H���  �҃�]�������������U��p3�H���   ��]������������U��EP�MQ�p3�B��l  �у�]����������������U��EP�p3�Q��   �Ѓ�]����U��EP�MQ�UR�p3�H��  �҃�]�������������U����M������E�P�p3�Q���   �Ѓ��M�Q�M������M�������E��]����������������U��p3�H��`  ��]������������U��EP�p3�Q��  �Ѓ�]����U����EP�M�Q�p3�B���   �у��U��
�H�J�H�J�H�J�H�J�@�B�E��]���U��EP�MQ�p3�B���  �у�]����������������U��EP���E�$���E�$�MQ�p3�B���   �у�]��������������U��EP�MQ�UR�p3�H���   �҃�]�������������U��EP�MQ�UR�p3�H���   �҃�]�������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�UR�p3�H���   �҃�]�������������U��EP�MQ�p3�B���   �у�]����������������U��EP�MQ�p3�B���   �у�]����������������U��EP�p3�Q���   �Ѓ�]����U��EP�p3�Q���   �Ѓ�]����U��EP�p3�Q���   �Ѓ�]����U����M��E�P�M�Q�U�R�E�P�p3�Q���   �Ѓ���u3���E��]�����U����M��E�P�M�Q�U�R�E�P�p3�Q���   �Ѓ���u3���E���]�����U����M��E�P�M�Q�U�R�E�P�p3�Q���   �Ѓ���u3���E���]�����U��EP�p3�Q��8  �Ѓ�]����U��Q�M��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�1g��P�U�R�p3�H0���   �҃�(��]�$ ���U��Q�M��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�aG  P�U�R�p3�H0���   �҃�(��]�$ ���U��Q�M��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P�p3�Q0���   �Ѓ�(��]�$ �������U��Q�M��EP�MQ�UR�EP�M�Q�p3�B0���   �у���]� �����������U��Q�M��E�P�p3�Q0���   �Ѓ���]��������������U��Q�M��EP�MQ�U�R�p3�H0���   �҃���]� ����U��Q�M��EP�MQ�UR�EP�M�Q�p3�B0���   �у���]� �����������U��Q�M��E�P�p3�Q0���   �Ѓ���]��������������U��p3�H0���   ��]������������U��E�Q�p3�B0���   �у��U�    ]���������U��EP�p3�Q��H  �Ѓ�]����U��EP�p3�Q��T  �Ѓ�]����U��p3�H��p  ��]������������U��p3�H���  ��]������������U��EP�p3�Q���  �Ѓ�]����U��EP�p3�Q���  �Ѓ�]����U��EP�p3�Q���  �Ѓ�]����U��EP�MQ�UR�EP�p3�Q���  �Ѓ�]��������U��EP�MQ�UR�EP�MQ�p3�B���  �у�]����U����EP�MQ�UR�E�P�p3�Q��X  �Ѓ�P�M�m����M������E��]���������������U���$j hLGOg�M������PhicMC�E�P�������M������M�艫����u�M�m����M������E��M��h���P�M�����M������E��]�U��EP�MQ�p3�B��  �у�]����������������U��EP�p3�Q��\  �Ѓ�]����U����EP�MQ�U�R�p3�H��t  �҃����o���M��n���E��]������U����EP�M�Q�p3�B���  �у�P�M蕑���M�轏���E��]�������U����EP�M�Q�p3�B���  �у�P�M�U����M��}����E��]�������U��EP�p3�Q���  �Ѓ�]����U��EP�p3�Q���  �Ѓ�]����U��EP�p3�Q���  �Ѓ�]����U��E$P�M Q�UR�EP�MQ�UR�EP�MQ�p3�B���  �у� ]��������U��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�p3�H���  �҃�$]�����U���j �EP�MQ�UR�EP�M�Q�p3�B��t  �у�P�M�'����M��O����E��]���������U����EP�MQ�UR�EP�M�Q�p3�B���  �у�P�M�i����M������E��]�����������U��EP�p3�Q��8  �Ѓ�]����U���  �p!3ŉE��E�E��M�Q�URh   ������P�	  ��������Qhh��p3�B��4  �у��E�    �M�3��k�  ��]�������U����E�P�p3�Q��  �Ѓ�P�M�	����M��1����E��]�����������U����E�P�p3�Q��  �Ѓ�P�M�Ɏ���M������E��]�����������U���(������u�Vh���M������EPh���M��q����MQh���M��`���j �U�RhicMC�E�P�L������M������M��������]������U���(�%�����u�M�	����E�Xh!���M��7����EPh!���M������j �M�QhicMC�U�R����������h���P�M�ߍ���M������M��O����E��]���������U���(������u�M艍���E�Xh����M������EPh����M��v���j �M�QhicMC�U�R�b�����������P�M�_����M������M�������E��]���������U���(�%�����u3��Rh#���M��@����EPh#���M������j �M�QhicMC�U�R����������Q����E�M������M��^����E��]��������U���(������u3��Rhs���M�������EPhs���M�菍��j �M�QhicMC�U�R�{�������������E�M������M�������E��]��������U��EP�MQ�UR�EP�MQ�UR�p3�H���  �҃�]�U��EP�MQ�UR�p3�H��@  �҃�]�������������U��EP�MQ�UR�EP�MQ�UR�p3�H���  �҃�]�U��E�8 t�M�R�p3�H��D  �҃��E�     ]��U��EP�p3�Q��H  �Ѓ�]����U��EP�p3�Q��L  �Ѓ�]����U��EP�MQ�UR�p3�H��P  �҃�]�������������U��EP�MQ�UR�p3�H��T  �҃�]�������������U��EP�MQ�UR�p3�H��X  �҃�]�������������U��EP�MQ�UR�p3�H��\  �҃�]�������������U��p3�H��d  ��]������������U��E P�MQ�UR�EP�MQ�UR�EP�p3�Q��h  �Ѓ�]������������U��EP�MQ�p3�B��l  �у�]����������������U��p3�H���  ��]������������U����EP�M�Q�p3�B���  �у�P�M�����M��=����E��]�������U��EP�p3�Q���  �Ѓ�]����U��EP�p3�Q���  �Ѓ�]����U��EP�MQ�p3�B���  �у�]����������������U��EP�p3�Q���  �Ѓ�]����U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�MQ�UR�p3�H��l  �҃�]�������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��EP�p3�Q���  �Ѓ�]����U��EP�MQ�p3�B��$  �у�]����������������U��EP�p3�Q��(  �Ѓ�]����U��EP�p3�Q��,  �Ѓ�]����U��p3�H��0  ��]������������U��p3�H��<  ��]������������U��EP�MQ�UR�EP�p3�Q���  �Ѓ�]��������U��p3�H���  ��]������������U��EP�MQ�UR�p3�H���  �҃�]�������������U��]������������U��E$P�M Q�UR�EP�MQ�UR�EP�MQ�p3�B��  �у� ]��������U��p3�H��P  ��]������������U��EP�MQ�UR�p3�H��`  �҃�]�������������U��Q�M��E���P�}   ����]�������U��Q�} 3��Z�EP�MQ�UR�EP覲  ���E��}� |�M��9M�|+�}� }hp�hH  �q������UU�B� �E���E��E���]�����U��EP�p3���   ���   �Ѓ�]�U��EP�MQ�p3�Bd�HP�у�]���U��E�8 u��MQ�p3�Bd�HT�у�]�������������U��Q�M��EP�MQ�UR�EP�M�Q�p3�Bh��у���]� ���������������U��Q�M��EP�MQ�UR�EP�M�Q�p3�Bh���   �у���]� �����������U��Q�M��EP�MQ�UR�E�P�p3�Qh�B�Ѓ���]� ��U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�Hh�Q �҃���]� �����������U��Q�M��EP�MQ�UR�EP�M�Q�p3�Bh���   �у���]� �����������U��Q�M��EP�M�Q�p3�Bh���   �у���]� �������U��p3�Hh�QX��]���������������U��E�8 u��MQ�p3�Bh�H\�у�]�������������U��Q�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�p3�Bh�H`�у� ��]� ��U��Q�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�p3�Bh�Hd�у� ��]� ��U��Q�M��EP�MQ�U�R�p3�Hh�Qh�҃���]� �������U��Q�M��EP�MQ�U�R�p3�Hh�Ql�҃���]� �������U��Q�M��EP�MQ�U�R�p3�Hh�Qp�҃���]� �������U��Q�M��EP�MQ�UR�E�P�p3�Qh�Bt�Ѓ���]� ��U��EP�MQ�UR�EP�MQ�p3�Bh���   �у�]����U��Q�M��EP�M�Q�p3�Bh�Hx�у���]� ����������U��Q�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�p3�Bh���   �у� ��]� ���������������U��Q�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�p3�Bh���   �у� ��]� ���������������U��Q�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�p3�Bh���   �у� ��]� ���������������U��Q�M��EP�MQ�UR�E�P�p3�Qh�B|�Ѓ���]� �U��Q�M��E P���E�$���E�$���E�$�M�Q�p3�Bh���   �у� ��]� ������������U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�Hh���   �҃���]� ��������U��Q�M��EP�MQ�UR�EP�M�Q�p3�Bh���   �у���]� �����������U��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�p3�Hh���   �҃�$]�����U��E<P�M8Q�U4R�E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�p3�Bh���   �у�8]����������������U��E@P�M<Q�U8R�E4P�M0Q�U,R�E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�p3�Hh���   �҃�<]�������������U���(�M؍M���V���EP�M�����P�M��Z���j �M�Q�U�R�M��x����M�������E�P�M�t����M������E��]� ���U��Q�M��EP���E�$�M�Q�p3�Bh���   �у���]� ��������������U��Q�M��EP���E�$�M�Q�p3�Bh���   �у���]� ��������������U��Q�M��EP�MQ�U�R�p3�Hh���   �҃���]� ����U��Q�M��EP�MQ�U�R�p3�Hh���   �҃���]� ����U����M�E(P�M$Q���E�$���E�$�UR�EP�M�Q�U�R�p3�Hh���   �҃�(�M���P�Q�P�Q�P�Q�P�Q�@�A�E��]�$ ������������U����M�E$P���E�$���E�$�MQ�UR�E�P�M�Q�p3�Bh���   �у�$�U��
�H�J�H�J�H�J�H�J�@�B�E��]�  ���������������U��p3�HL���   ��]������������U��E�Q�p3�B@�H�у��U�    ]������������U��p3�HL���]����������������U��E�Q�p3�B@�H�у��U�    ]������������U��Q�M��E�P�p3�QL���   �Ѓ���]��������������U��Q�M��EP�MQ�U�R�p3�HL���   �҃���]� ����U����M��E�P�p3�QL���   �Ѓ��E��}� uj �MQ�U�R�p3�HL���   �҃���M��?   P�M�������]� U��Q�M��E�P�p3�QL��(  �Ѓ���]��������������U��Q�M��EP�MQ�U�R�p3�HL��,  �҃���]� ����U��p3�HL�Q��]���������������U��E�Q�p3�B@�H�у��U�    ]������������U����M�EP�M�Q�U�R�p3�HL�Q�҃�P�M�����M��*����E��]� �U��Q�M��EP�M�Q�p3�BL���   �у���]� �������U��Q�M��EP�MQ�U�R�p3�HL�Q�҃���]� �������U��Q�M��E�P�p3�QL�B�Ѓ���]�U��Q�M��E�P�p3�QL�B�Ѓ���]�U��Q�M��E�P�p3�QL�B�Ѓ���]�U��Q�M��EP�MQ�UR�E�P�p3�QL�B �Ѓ���]� ��U��Q�M��EP�M�Q�p3�BL��4  �у���]� �������U��Q�M��EP�MQ�UR�E�P�p3�QL�B$�Ѓ���]� ��U��Q�M��EP�MQ�UR�EP�M�Q�p3�BL�H(�у���]� ��������������U��Q�M��E�P�p3�QL�B,�Ѓ���]�U��Q�M��E�P�p3�QL�B0�Ѓ���]�U��Q�M��EP�MQ�U�R�p3�HL��  �҃���]� ����U��Q�M��E�P�p3�QL���   �Ѓ���]��������������U����M�EP�M�Q�U�R�p3�HL��  �҃�P�M�����M������E��]� ��������������U��Q�M��E�P�p3�QL�B4�Ѓ���]�U��Q�M�j �E�P�p3�QL�B8�Ѓ���]���������������U��Q�M��EP�MQ�p3�BL�M����   �ҋ�]� �������U��Q�M��EP�MQ�p3�BL�M����   �ҋ�]� �������U��Q�M��EP�MQ�p3�BL�M����   �ҋ�]� �������U��Q�M��EP�MQ�p3�BL�M����   �ҋ�]� �������U��Q�M��EP�MQ�p3�BL�M����   �ҋ�]� �������U��Q�M��EP�MQ�p3�BL�M����   �ҋ�]� �������U��Q�M��EP�MQ�UR�EP�p3�QL�M���l  �Ћ�]� ���������������U��Q�M��EP�p3�QL�M����   �Ћ�]� �����������U��Q�M��EP�p3�QL�M����   �Ћ�]� �����������U��Q�M��EP�p3�QL�M����   �Ћ�]� �����������U��Q�M��EP�M�Q�p3�BL�H<�у���]� ����������U��Q�M��E�P�p3�QL�B�Ѓ���]�U��Q�M��EP�MQ�U�R�p3�HL�Q@�҃���]� �������U��Q�M�j �EP�M�Q�p3�BL�HD�у���]� ��������U��Q�M�j �EP�M�Q�p3�BL�HH�у���]� ��������U��Q�M�j�EP�M�Q�p3�BL�HD�у���]� ��������U��Q�M�j�EP�M�Q�p3�BL�HH�у���]� ��������U���4�M̍M��oL��h�  �M�����P�M��ɷ��j �E�P�M�Q�M�����������E�M��%����U��t�E�    �M��n����E���M������EЍM��V����EЋ�]����������������U���(�M�j�M��E��h�  �M�����P�M��7���j�E�P�M�Q�M�腓���M�蝸���M��������]��U���(�M؋EP�M��k  h�  �M��.���P�M�����j�M�Q�U�R�M��3����M��K����M�������]� �������������U���(�M؋EP�M��  h�  �M������P�M�腶��j�M�Q�U�R�M��Ӓ���M������M��C�����]� �������������U���,�MԍM���J��h�  �M��r���P�M��)���j �E�P�M�Q�M��G���������E�M�腷���U��t�M�eN���M�������E��M��  P�M�O���M������E��]� ������U���,�MԍM��?J��h�  �M������P�M�虵��j �E�P�M�Q�M�跑��������E�M�������U��t�M��M���M��=����E��M��   P�M�N���M������E��]� ������U���<�MčM��I��h�  �M��R���P�M��	���j �E�P�M�Q�M��'���������E�M��e����U��t���]ЍM������E���M��  �]ȍM������Eȋ�]��U���4�M̍M��/I��h�  �M������P�M�艴��j �E�P�M�Q�M�觐��������E�M������U��t�E�    �M��.����E���M��Q����EЍM������EЋ�]����������������U���,�MԍM��H��h�  �M��B���P�M������j �E�P�M�Q�M�����������E�M��U����U��t�M�C���M������E�,�M���  �M���P�Q�P�Q�@�A�M��o����E��]� ������U��Q�M��E�P�p3�QL���   �Ѓ���]��������������U����M�j�EP�M�Q�U�R�p3�HL���   �҃��M���P�Q�P�Q�@�A�E��]� ����U����M�j �EP�M�Q�U�R�p3�HL���   �҃��M���P�Q�P�Q�@�A�E��]� ����U���,�MԍM��/G��h�  �M������P�M�色��j �E�P�M�Q�M�觎��������E�M������U��t�M�%B���M��-����E�,�M��P  �M���P�Q�P�Q�@�A�M�������E��]� ������U���,�MԍM��F��h�  �M��2���P�M�����j �E�P�M�Q�M�����������E�M��E����U��t�M�A���M������E�,�M��  �M���P�Q�P�Q�@�A�M��_����E��]� ������U���,�MԍM���E��h�  �M�����P�M��I���j �E�P�M�Q�M��g���������E�M�襲���U��t�M��@���M�������E�,�M��  �M���P�Q�P�Q�@�A�M������E��]� ������U���4�M̍M��OE��h�  �M������P�M�詰��j �E�P�M�Q�M��ǌ��������E�M������U��t�E�    �M��N����E���M��q����EЍM��6����EЋ�]����������������U���(�M؃��E�$�M��f  h�  �M��Y���P�M�����j�E�P�M�Q�M��^����M��v����M��������]� ��������U���(�M؋EP�M��=��h�  �M������P�M�赯��j�M�Q�U�R�M������M������M��s�����]� �������������U���(�M؋EP�M���  h�  �M�螿��P�M��U���j�M�Q�U�R�M�裋���M�軰���M�������]� �������������U���(�M؋EP�M��{  h�  �M��>���P�M������j�M�Q�U�R�M��C����M��[����M�������]� �������������U���(�M؋EP�M��  h�  �M��޾��P�M�蕮��j�M�Q�U�R�M������M�������M��S�����]� �������������U���(�M؋EP�M��  h�  �M��~���P�M��5���j�M�Q�U�R�M�胊���M�蛯���M��������]� �������������U���(�M؋EP�M��;��h�  �M�����P�M��խ��j�M�Q�U�R�M��#����M��;����M�������]� �������������U���,�MԍM��B��h�  �M��½��P�M��y���j �E�P�M�Q�M�藉��������E�M��ծ���U��t�M�=���M������E�,�M��@  �M���P�Q�P�Q�@�A�M�������E��]� ������U���4�M̍M��A��h�  �M��"���P�M��٬��j �E�P�M�Q�M������������E�M��5����U��t�E�    �M��~����E���M������EЍM��f����EЋ�]����������������U���4�M̍M���@��h�  �M�蒼��P�M��I���j �E�P�M�Q�M��g���������E�M�襭���U��t�E�    �M�������E���M������EЍM�������EЋ�]����������������U����M��M�������E��}�t�}�t�}�t	�E�    ��E�   �E��]����U��Q�M��p3�PL�M����  �Ћ�]���U���(�M؋EP�M���  h�  �M�螻��P�M��U���j�M�Q�U�R�M�裇���M�軬���M�������]� �������������U���(�M؋EP�M���8��h�  �M��>���P�M������j�M�Q�U�R�M��C����M��[����M�������]� �������������U���(�M؋EP�M��k8��h�  �M��޺��P�M�蕪��h�   j�I<����P�M�Q�U�R�M��Ն���M������M��E�����]� ���������������U��EP�p3�Q���   �Ѓ�]����U��EP�p3�Q���   �Ѓ�]����U��p3�H���   ��]������������U��p3�H���   ��]������������U��E�Q�p3�B���   �у��U�    ]���������U��EP�p3�Q���   �Ѓ�]����U��Q������E��}� u3��Oj �EP�MQ�UR�E�P�p3�Q��h  �Ѓ���u"�}� t�M�Q�p3�B@�H�у��E�    �E���]��������U��j �EPj �MQ�:����P�UR�EP�p3�Q��h  �Ѓ�]�����������U��EP�MQ�UR�EP�p3�Q���   �Ѓ�]��������U��E P�MQ�UR�EP�MQ�UR�EP�p3�Q���   �Ѓ�]������������U��Q�M��E�P�p3�QL�BL�Ѓ���]�U��Q�M��E�P�p3�QL�BP�Ѓ���]�U��Q�M��EP�MQ�UR�E�P�p3�QL���  �Ѓ���]� ���������������U��Q�M��EP�M�Q�p3�BL��  �у���]� �������U��Q�M��EP�M�Q�p3�BL���   �у���]� �������U��Q�M��E�P�p3�QL�BX�Ѓ���]�U��Q�M��EP�MQ�UR�E�P�p3�QL�B\�Ѓ���]� ��U���L�M������E��}� u3��^  �E�    �E�    �E�    �M�蕺���M��	  �E��E܍MȉM�URh]  �M��@5��j j �E�P�M���	  ��u�   �M������E���MĉM��}� ��   �M��"����EċU��U��E�Ph�   ��������u�w�}� u�oj �M��	  �E��}� u�Z�M�Q�M��	  �U�R�������}� t�E�P�p3�Q@�B�Ѓ��E�    �l����M��M��M��H����M��0����E��G�}� t�U�R�p3�H@�Q�҃��E�    �E�P�������E�    �M�������M������E���]� ��������������U��Q�M��E�P�p3�QL�B`�Ѓ���]�U��Q�M��E�P�p3�QL�Bd�Ѓ���]�U��Q�M��EP�M�Q�p3�BL�Hh�у���]� ����������U��Q�M��E�P�p3�QL��D  �Ѓ���]��������������U��Q�M��E�P�p3�QL�Bl�Ѓ���]�U��Q�M��EP�M�Q�p3�BL���   �у���]� �������U��Q�M��E��M�H�U��E$�Bhбh��h��hp��M��QR�E P�MQ�UR���E�$�EP�M��QR�E�P�p3�QL���   �Ѓ�4��]�  ��������������U��E��M���]����������������U��EP�M��M�B��]�����������U��EP�MQ�U��M�P��]�������U��EP�MQ�UR�EP�M��M�B��]���������������U��Q�M��E�P�p3�QL���   �Ѓ���]��������������U��Q�M��EP�MQ�UR�E�P�p3�QL��   �Ѓ���]� ���������������U��Q�M��EP�MQ�UR�EP�MQ�p3�BL�M���H  �ҋ�]� �����������U��Q�M��p3�PL�M���L  �Ћ�]���U��Q�M��EP�p3�QL�M���P  �Ћ�]� �����������U��Q�M��EP�p3�QL�M���T  �Ћ�]� �����������U��Q�M��EP�MQ�p3�BL�M���p  �ҋ�]� �������U��Q�M��EP�MQ�p3�BL�M���t  �ҋ�]� �������U��Q�M��EP�MQ�UR�EP�MQ�U�R�p3�HL���   �҃���]� ��������U��Q�M��EP�MQ�UR�E�P�p3�QL���   �Ѓ���]� ���������������U��Q�M��EP�MQ�UR�EP�M�Q�p3�BL��   �у���]� �����������U���(�M���  �M���  �} t�M��,  ��u�E�   �M���  �M��Q����E��Kj�M��  P�M�����M���  �E��E�E�M�Qh=����������E؍M��  �M������E؋�]��������������U���(�M��R  �M��:  �} t�M��  ��u�E�   �M��Y  �M������E��Kj�M��b  P�M������M��Q  �E��E�E�M�Qh<���Z������E؍M��  �M��d����E؋�]��������������U��EP�MQ�UR�p3�HL���   �҃�]�������������U��EP�MQ�p3�BL���   �у�]����������������U��EP�MQ�p3�BL���   �у�]����������������U��p3�HL��  ��]������������U��p3�HL��@  ��]������������U��Q�M��EP�MQ�p3�BL�M����  �ҋ�]� �������U��Q�M��EP�MQ�p3�BL�M����  �ҋ�]� �������U��Q�M��EP�p3�QL�M����  �Ћ�]� �����������U��Q�M��p3���   �M��BP�Ћ�]���U��Q�M��E��     �M��A    �UR�E�P�p3���   �B(�Ѓ��E���]� �U��Q�M��E�P�p3���   �BL�Ѓ���]��������������U��Q�M��E�P�p3���   �B<�Ѓ���]��������������U��Q�M��E�P�p3���   �BP�Ѓ���]��������������U��Q�M��E��    �M��E�Y�E���]� ��������������U��Q�M��E��     �M��A    �UR�E�P�p3���   �B,�Ѓ��E���]� �U��Q�M��E��     �M��A    �U��B    �E��@    �M��A    �U��B    �E��@    �E���]��������������U��Q�M��EP�MQ�UR�p3���   �M��B�Ћ�]� ����U��Q�M��EP�p3���   �M����   �Ћ�]� ��������U��Q�M��EP�p3���   �M��B<�Ћ�]� �����������U��Q�M��   �M���E���]���������U��p3���   ���   ��]���������U��Q�M��E�P��������M��    ��]�U��Q�M��E�� ��]�U��Q�M��h��]����z	�h��]�`��]����Au	�`��]�E���X����$�+�����E���M����Y�M���  �E���]� ��������U����M����]����Az	�E�   ��E�    ���]����Az	�E�   ��E�    �E�3�;E����M����E�$�C  ���X����$�*�����U�����E�$�  ���X����$�U*�����E��X�M����Y����Auh��j��������U����Z�}� u�E�� ���M���M���   �E���]� ���U��Q�M��E��E�X�M����Y����Auh�j,�u������U����Z��]� ����U����M����]����Auh0�j5�?��������]�E�� �M���$�)�����M����A�$�]��m)�����}���$�\)�����U�����E�$�F)�����E��X�M��   ��]� ���������������U���4�M̋Ẽ�� �$�  ���]��M̃��A�$�  ���]��P��]�����At�P��]�����Au�U�����E����X�U  �x��]�����Auz�x��]�����Auj�E���:  �E��E���:  �E��}� u�M�����U����Z�8�Eܙ�}��U�E��E܋M�M��}� u��E܋U��:�E���E܋M��y�U��Z��   ���E��$���E��$��   ���=p��]����]�����Au.�E��M��]��E��M��]��E�� �MЋM���U��B�MЋE��X���]�����Au���]��M����Y���E��$���E��$�   ���]��E��]��E��]��X��]�����A{ǋU���u��E���M��A�u��U��Z��]��������������U����E�$�J  ��]�����������U���E�]����Au�E��E]�������U����E�$���E�$�&K  ��]��U��E��M�B��]���������������U��E��M�B��]���������������U��Q�M��E�� ���M��A    h���U�RhP�h0��p3�HP��҃��M��A�E���]��������U��E��M�B��]���������������U��Q�M��E�� ���M��y u�U��BP�p3�QP�B�Ѓ���]������������U��Q�M��E��x u3��"j �MQ�UR�E��HQ�p3�BP�H�у���]� ����U��Q�M��E��x t�MQ�U��BP�p3�QP�B�Ѓ���]� ��������������U��Q�M��E��x t�MQ�U��BP�p3�QP�B�Ѓ���]� ��������������U��p3�HP���   ��]������������U��EP�p3�QP���   �Ѓ�]����U��p3�HP�QP��]���������������U��EP�p3�QP�BT�Ѓ�]�������U��Q�M��E��     �M��A    �E���]����������������U��Q�M��E��8 u�6�M��R�p3�HP�QL�҃��E��Q�p3�BP�H<�у��U��    ��]������U��Q�M��EP�MQ�M�  P�M��   ��]� ����������U����M��E��8 t)�M��R�p3�HP�Q<�҃��E��     �M��A    �U��E�Bh���MQhP�h0��UR�EP�p3�QP�B8�Ѓ��M���E�    �	�U����U��E�;E}f�M��U���x u.�M��U���@   �M��U���HQ�p3�BP�H�у��U�R�E��Q�p3�BP�H@�у��U��M���B뉋E�3Ƀ8 ������]� ���������U����M��E�    �E�    �	�E����E��M�U�;Q}a�E�P�M�R�p3�HP�Q@�҃��E��}� t!j �EPj�M�Q�p3�BP�H�у���u�U�P�p3�QP�BL�Ѓ�3��닸   ��]� �������U��Q�M��E��Q�p3�BP�HD�у���]���������������U��Q�M��E��Q�p3�BP�HH�у���]���������������U��Q�M��E��Q�p3�BP�HL�у���]���������������U��Q�M�3���]����U��Q�M��M��q����E��t�M�Q�`�����E���]� ����U��Q�M��E��@��]����������������U��Q�E�E��}�t��M��3�U��3�   ��]� �U����E�E��M����M��}��>  �U��$�D��   �-  ��3����3�=�3��   �MQ��g����=�6  }
�������   �} u
�������   h��jmh�3j�S�����E��}� t�M��)���E���E�    �U��3�=�3 t�EP��3��-���   �   �MQ�UR�KK������u����o�   �h�#K���a��3����3uH�=K���h\���=�3 t+��3�M�U�U��}� tj�M�� e���E���E�    ��3    �   ������]������	�=�������U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U����M�E�P�M�Q�p3�BX��у��U��
�H�J�H�J�H�J�H�J�@�B�E��]� �U����M�E�P�M�Q�p3�BX�H�у��U��
�H�J�H�J�H�J�H�J�@�B�E��]� U����M�E�P�M�Q�p3�BX�H�у��U��
�H�J�H�J�H�J�H�J�@�B�E��]� U���dVW�M��E�P�M�Q�p3�BX�H�у��   ���}�E_^��]� �����U��Q�M��EP�M�Q�p3�BX�H�у���]� ����������U��Q�M��EP�M�Q�p3�BX�H�у���]� ����������U��Q�M��EP�M�Q�p3�BX�H�у���]� ����������U��Q�M��EP�M�Q�p3�BX�H�у���]� ����������U��Q�M��EP�M�Q�p3�BX�H$�у���]� ����������U��Q�M��EP�M�Q�p3�BX�H �у���]� ����������U��Q�M��EP�MQ�U�R�p3�HD�Q�҃���]� �������U��j �EP�p3�QD��Ѓ�]������U��E�Q�p3�B@�H�у��U�    ]������������U��EP�MQ�p3�BD��у�]����U��E�Q�p3�B@�H�у��U�    ]������������U��j �EP�p3�QD��Ѓ�]������U��E�Q�p3�B@�H�у��U�    ]������������U��EPh2  �p3�QD��Ѓ�]���U��E�Q�p3�B@�H�у��U�    ]������������U��EPhO  �p3�QD��Ѓ�]���U��E�Q�p3�B@�H�у��U�    ]������������U��EPh'  �p3�QD��Ѓ�]���U��E�Q�p3�B@�H�у��U�    ]������������U��j h�  �p3�HD��҃�]������U��E�Q�p3�B@�H�у��U�    ]������������U��j h:  �p3�HD��҃�]������U��E�Q�p3�B@�H�у��U�    ]������������U����M�M��  �E�    �E�    �E�Pj�M��C�����u3���E���]�����U��j h�F �p3�HD��҃�]������U��E�Q�p3�B@�H�у��U�    ]������������U��j h�_ �p3�HD��҃�]������U��E�Q�p3�B@�H�у��U�    ]������������U����M�} u3��0�M��  �E�    �E�E��M�Qj�M��Z����u3���   ��]� �������U��Q�M��E�P�p3�QD�B$�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E�P�p3�QD�B(�Ѓ���]�U��Q�M��E�P�p3�QD�B�Ѓ���]�U��Q�M��E��     �M��A    �E���]����������������U��Q�M��E��     �M��A    �U��B    �E��@    �E���]������������U��Q�M��M��1  ��]��������������U��Q�M��E��     �M��A    �U��B    �E��@    �M�U�A;BuKjj�M��  ��u�   �M���E��
�U���M�Q�P�E���U�B�A�M��Q�   �Tjj�M���   ��u�B�E���U���M���E�H�J�U���M�Q�P�E���U�B�A�M��Q�   �E���]� ������������U��Q�M��E��     �M��A    �U��B    �E��@    �MQ�M��6  �E���]� �������������U��Q�M��EP�M��  �E���]� ����U��Q�M��M��   �} ��   h��jI�E��P�p3�Q���   �Ѓ��M���U��: u3��b�} tAh��jN�E��P�p3�Q���   �Ѓ��M��A�U��z u�E�P�o����3���M��U�Q�E��M�H�   �3���]� ������������U��Q�M��E�P��n�����M���Q�n�����U��B    �E��@    ��]�������U��Q�M��M������} ��   �E�8 ��   �M�y ��   h�jl�U�B��P�p3�Q���  �Ѓ��M���U��: u3��   �E�x tI�M�y t@h<�jq�U�B��P�p3�Q���  �Ѓ��M��A�U��z u�M�����3��^�E��M�Q�P�E��M�Q�P�E��HQ�U��P�M�R�  ���E��x t�M��QR�E��HQ�U�BP�m  ���   ��]� ���������������U��Q�M��M������} �9  �} �/  hh�h�   �E��P�p3�Q���  �Ѓ��M���U��: u3���   �} tT�} tNh��h�   �E��P�p3�Q���  �Ѓ��M��A�U��z u�M������3��   �E��M�H�M�U��B   h��h�   �E��H��Q�p3�B���  �у��U��B�E��x u�M�����3��T�M��U�Q�E��HQ�U��P�MQ�.  ���} t�U��BP�M��QR�EP�  ����M��Q�E��   ��]� ���U��Q�M��E��     �M��A    �U��B    �E��@    ��]���������������U���  VW��|������]��E�    j �M�艈��j �M�����j �M��u�����|����H�U�<�}���]  �} ��  �M��=��j ��x����=�����|�����k�U��EȋJ�M̋B�EЋJ�MԋB�E؋J�M܍U�R��|�����Qk�UR��`���P舁�������x����P��|����H�M��P�U��H�M��P�U��E�   �	�E����E���|����Q�E�;��   �M�Q��|�����M���k�UR��H���P��������M��P�U��H�M��P�U��H�M��P�UčE�P��x���Q��0���R�~����P�M��h  �E���x����M���|����U��U��E��E��M��M��UĉU��F��������$����������E������������P�� ����H��$����P��(����H��,����P�E�P�� ���Q��~�����U��H��
�H�J�H�J�H�J�H�J�@�B���E��$�u����E��$ݝt����d�����ܝt���������   ���E��$�B����E��$ݝl����1�����ܝl���������   �M��HQ�����$�����$�����$�������3;��P������R�6}�����M�����P�Q�P�Q�P�Q�P�Q�@�A�M��Q�U��HR������P��|�����M��0���P�Q�P�Q�P�Q�P�Q�@�A�  ���E��$�c����E��$ݝd����R�����ܝd���������   �����$�����$�����$�������[:��P�M��HQ������R�W|�����M�����P�Q�P�Q�P�Q�P�Q�@�A�M��Q�U��HR��p���P�|�����M��0���P�Q�P�Q�P�Q�P�Q�@�A�   �����$�����$�����$��X����9��P�M��HQ��@���R�{�����M��0���P�Q�P�Q�P�Q�P�Q�@�A�M��HQ�U��0R��(���P�f{�����M�����P�Q�P�Q�P�Q�P�Q�@�A�MQ������R������   ���}��E�    �	�E����E��M�;M}��|����B�M��U���U��؋�|�����U���k�EP�MQ������R��  ����MȋP�ŰH�MЋP�UԋH�M؋P�U܋�|�����U��D�k�EP�MQ������R�  ����M��P�U��H�M��P�U��H�M��P�U��E�    �	�E����E���|����Q�E�M�;���   �E�����|����J�u��<�U���|������k�UR�EP������Q�  ����U�H�M�P�U��H�M�P�U��@�E��M�Q�U�R�E�P�h   ���E��]��M��MȋU��ŰE��EЋM��MԋU��U؋EĉE܋M�M��U�U��E��E��M�M��U��U��E��E������E�_^��]� �������U��E�M�@�a�U�
�E�M�@�a�U�
���E�M�@�a�U�
��]�����U��Qj�%   ���E��}� u3���E��H�ы�]����������U��h�3�EPh_� �
  ��]������U����E�8 u�5j��������E��}� u� �M��U��E�P�M��Q�҃��E�     ��]��������U����M�j�������E��}� t	�E��x u3���MQ�U��M��B�Ћ�]� ��U����M�j�@������E��}� t	�E��x u3���MQ�U��M��B�Ћ�]� ��U����M�j� ������E��}� t	�E��x u3���MQ�UR�EP�U��M��B�Ћ�]� ����������U����M�j�������E��}� t	�E��x u3���MQ�U��M��B�Ћ�]� ��U����M�j �p������E��}� t	�E��x  u3���MQ�U��M��B �Ћ�]� ��U����M�j$�0������E��}� t	�E��x$ u2���MQ�U��M��B$�Ћ�]� ��U����M�j(��������E��}� t	�E��x( u3���U��M��B(�Ћ�]���������U����M�j,�������E��}� t	�E��x, u3���U��M��B,�Ћ�]���������U����M�j0�p������E��}� t	�E��x0 u3���MQ�U��M��B0�Ћ�]� ��U����M�j4�0������E��}� t	�E��x4 u�����MQ�UR�E��M��P4�ҋ�]� �������������U����M�j8��������E��}� t	�E��x8 u3���U��M��B8�Ћ�]���������U����M�j<�������E��}� t	�E��x< u��MQ�U��M��B<�Ћ�]� ����U����M�j@�`������E��}� t	�E��x@ u��MQ�U��M��B@�Ћ�]� ����U����M�jD� ������E��}� t	�E��xD u3���MQ�U��M��BD�Ћ�]� ��U����M�jH��������E��}� t	�E��xH u��MQ�U��M��BH�Ћ�]� ����U����M�jL�������E��}� t	�E��xL u3���U��M��BL�Ћ�]���������U����M�jP�`������E��}� t	�E��xP u3���U��M��BP�Ћ�]���������U����M�jT� ������E��}� t	�E��xT u��U��M��BT�Ћ�]�����������U����M�jX��������E��}� t	�E��xX u��U��M��BX�Ћ�]�����������U����M�j\�������E��}� t	�E��x\ u��U��M��B\�Ћ�]�����������U����M�j`�`������E��}� t	�E��x` u3���MQ�UR�E��M��P`�ҋ�]� ��������������U����M�jd�������E��}� t	�E��xd u3���MQ�UR�E��M��Pd�ҋ�]� ��������������U����M�jh��������E��}� t	�E��xh u��MQ�UR�EP�MQ�UR�E��M��Ph�ҋ�]� ����U����M�jl�p������E��}� t	�E��xl u3���MQ�UR�EP�U��M��Bl�Ћ�]� ����������U����M�jp� ������E��}� t	�E��xp u3���MQ�UR�E��M��Pp�ҋ�]� ��������������U����M�jt��������E��}� t	�E��xt u3���MQ�UR�E��M��Pt�ҋ�]� ��������������U����M�jx�������E��}� t	�E��xx u3���MQ�UR�E��M��Px�ҋ�]� ��������������U����M�j|�0������E��}� t	�E��x| u3���MQ�U��M��B|�Ћ�]� ��U����M�h�   ��������E��}� t�E����    u3���MQ�UR�E��M����   �ҋ�]� �����U����M�h�   �������E��}� t�E����    u����&�MQ�UR�EP�MQ�UR�EP�U��M����   �Ћ�]� ����U����M�h�   �=������E��}� t�E����    u����&�MQ�UR�EP�MQ�UR�EP�U��M����   �Ћ�]� ����U����M�h�   ��������E��}� t�E����    u3���MQ�UR�EP�MQ�U��M����   �Ћ�]� �������������U����M�h�   �}������E��}� t�E����    u3���MQ�U��M����   �Ћ�]� ���������U����M�h�   �-������E��}� t�E����    u��MQ�U��M����   �Ћ�]� �����������U����M�h�   ��������E��}� t�E����    u3���MQ�UR�E��M����   �ҋ�]� �����U����M�h�   �������E��}� t�E����    u3���MQ�UR�EP�U��M����   �Ћ�]� �U���   ��L����M���+���E�    �	�E���E䋍L����U�;Q�  ��L�����U���"b����u�̋�L�����U����a����E�E��E��M��P;Quc�E��k�MQ�U��Bk�EP�M�Q��o����P�U��k�EP�M��Qk�UR�E�P�o����P�M�Q�]m����P�M��1  �h�U��k�EP�M��Qk�UR�E�P�mo����P�M��Qk�UR�E��Hk�MQ��h���R�Co����P��P���P��l����P�M���  ������M�Q�UR�m�����E��]� ���������U���H�M��M��  �E�    �	�E����E��M��U�;Q��   �E���U����`����u�ҋE���U����h`����E�E��E��k�MQ�M���  �U��Bk�EP�M���  �M��Qk�UR�M��  �E��M��P;Qt�E��Hk�MQ�M��  �S����UR�EP�M��  ��]� ���U����M��E�    �E�x|�M�9 u3��?�E�    �	�U����U��E�M�;H}�U��M����  ��t	�U����U��͋E���]���������U����M��E�E��	�M����M��U��E�;B}!�M���E����K  ��t�E�+E����˃����]� �U����M��} |�E��8 u����<�E�    �	�M����M��U��E�;B}�M���E�����^��;Eu�E���Ѓ����]� ��U���S�M��E� �E�    �	�E����E��M�U�;Q}3�E��U����^��;Eu�]��E��U����  ��؈]���E���[��]� �����U����M��E�    �E�    �	�E����E��M�U�;Q} �E��U����s  ���t	�E����E��̋E���]�������������U����M��E�    �E�    �	�E����E��M�U�;Q}�E��U�����]����t	�E����E��͋E���]��������������U����M��E�    �	�E����E��M��U�;Q}�E���U���%����M���M������E�    �	�U����U��E��M�;H}}�U���M�����   �ue�E���U����]���E��E����E��	�M���M�U��E�;B}3�M���E����\��;E�u�M���E����   ��U���U����o�����]����������������U����M��M��\����E�E��M���  �E�E���E�}�wz�M��$�4��U�����E� ����\�M�U����M�U��B��E�M�U��B��M�U��B��-�M�U��B��M�U��B���M�U��B��M�U�����]� ����������������U����M�M��[���E��M��  �E��E;E�t	�}���u�M;M�t	�}���u�_�}���t�U�U��}���t�E�E��}��t�M��U����M���   �M���U�����   @�E���   �ыE���]� ��������U��Q�M��E��M� ��U���E��M�@�A�U��Z�E��M�@�A�U��Z�E���]� �������������U��E�M�@(�	�U�B�E�M�@@�I���U�E�BX�H�����$�M�U�A �
�E�@�M�U�A8�J���E�M�@P�I�����$�U�E�B��M��U�E�B0�H���M�U�AH�J�����$�M�$���E]���������U���4�M̋M���#���M̃���#��������$�M��pg���E̋M��U�P�M��H�U�P�M��H�U��P������$�M��6g���Ẽ��MЉ�UԉP�M؉H�U܉P�M��H�U�P�E��@0    �E̋�]�������������U��Q�M��E��x0 ��   �M�U�������Au
�E��M���U�E��@�Z����Au�M��U�B�Y�E�M��A�X����Au�U��E�@�Z�M�U��B�����z�E��M��X�U�E��@ �Z����z�M��U�B�Y �E�M��A(�X����z�U��E�@�Z(�`�M�U������A�B�A�B�A�B�A�B�I�J�U����E��
��J�H�J�H�J�H�J�H�R�P�E��@0   ��]� U���d�M��E��x0 ��   ���X��$�M���Q�U�R�E�P��e����P�M�Q��   ���U��
�H�J�H�J�H�J�H�J�@�B�MQ�U���R�E�P�f�����M���P�Q�P�Q�P�Q�P�Q�@�A�^�����$�M��e���M�U���E��A�U��Q�E��A�U��Q�E��A�M�U���A�B�A�B�A�B�A�B�I�J��]� ���U��E�@�M���$�M�A�M���$�U��M���$�M�� ���E]�����U��Q�M��E�� %    ��]������������U����M��M��   �E��}��u3��
�   �M�����]�����U��Q�M��E����   @t�����U��%���3ҹ   ���]���������������U��E��P�MQ�UR�I  ��]�����U��p3�H\���]����������������U��E�Q�p3�B\�H�у��U�    ]������������U��Q�M��E�P�p3�Q\�B�Ѓ���]�U��Q�M��E�P�p3�Q\�B�Ѓ���]�U��Q�M��EP�M�Q�p3�B\�H�у���]� ����������U��Q�M��EP�MQ�U�R�p3�H\�Q�҃���]� �������U��Q�M��EP�M�Q�p3�B\�H�у���]� ����������U��Q�M��E�P�p3�Q\�B�Ѓ���]�U��Q�M��EP�M�Q�p3�B\�H �у���]� ����������U��Q�M��EP�MQ�U�R�p3�H\�Q$�҃���]� �������U��Q�M��EP�MQ�UR�EP�M�Q�p3�B\�H`�у���]� ��������������U��Q�M��EP�M�Q�p3�B\�H0�у���]� ����������U��Q�M��EP�M�Q�p3�B\�H@�у���]� ����������U��Q�M��EP�M�Q�p3�B\�HD�у���]� ����������U��Q�M��EP�M�Q�p3�B\�HH�у���]� ����������U��Q�M��E�P�p3�Q\�B4�Ѓ���]�U��Q�M��EP�MQ�U�R�p3�H\�Q8�҃���]� �������U��Q�M��EP�M�Q�p3�B\�H<�у���]� ����������U����M�j �M�}���M��5����E�E�P�M�f���E�    �	�M����M��U�;U�}3�E�P�M�Qh����U�R�M��#����E�P�M�'���M�Q�M���뼋�]� ���U����M�E�P�M����}� |o�M��]����M�Q�M�q���}� tU�E�    �	�U���U�E�;E�};�M�Q�M�E���U�R�M�9���	�E����E��M�;M��U�R�M��j�����봸   ��]� �����������U��E�M��U�E�B�MQj�UR蝃����]���������U��   ]�������U����} t�E�8 t�M��Pj�UR躃�����E��}� u3��5�M�貄���E��}� u3�� �} t�E�M���U��E;B~3���E���]Ë�Q����  YË�U��V��������EtV��K��Y��^]� ����!��!���!s��!���!��!��!A��!1��!���!Ë�U�������} t�  ��]�������̃=�Q t-U�������$�,$�Ã=�Q t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$��jh��y-  �E��uz�6-  ��u3��8  �Z!  ��u�;-  ����,  ����Q�#,  ��3�P&  ��y�  ���N+  ��x ��(  ��xj �$  Y��u��3��   �\(  ��3�;�u[9=�3~���3�}�9=4u��%  9}u�,(  �  �,  �E������   �   3�9}u�=�!�t�v  ��j��uY�5  h  j�>"  YY��;�����V�5�!�5�3���Ѕ�tWV�n  YY� ���N��V�  Y�������uW�  Y3�@�i,  � jh��,  ����]3�@�E��u9�3��   �e� ;�t��u.�����tWVS�ЉE�}� ��   WVS�C����E����   WVS�����E��u$��u WPS����Wj S���������tWj S�Ѕ�t��u&WVS�������u!E�}� t�����tWVS�ЉE��E������E���E��	PQ�y.  YYËe��E�����3��q+  Ë�U��}u�t.  �u�M�U�����Y]� ��U��QSV�5�W�5�Q���5�Q�؉]��֋�;���   ��+��G��ruS�.  �؍GY;�sH�   ;�s���;�rP�u��   YY��u�C;�r>P�u��   YY��t/��P�4�����Q�u�=��׉��V�ף�Q�E�3�_^[�Ë�Vjj �   YY��V����Q��Q��ujX^Ã& 3�^�jh��*  �   �e� �u�����Y�E��E������	   �E��1*  ��   Ë�U���u���������YH]��������������̋T$�L$��ti3��D$��u���   r�=�Q t�-  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$Ë�U��S�]���woVW�=5 u��/  j�(.  h�   �  YY��t���3�@Pj �55������u&j^9L;tS�m0  Y��u���	0  �0�0  �0��_^�S�L0  Y��/  �    3�[]Ë�U��} t-�uj �55����uV�/  ����P�m/  Y�^]��������̃=�P ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�0  ��=�P t2���\$�D$%�  =�  u�<$f�$f��f���d$u��/  ���$��3  �   ��ÍT$�m3  R��<$tPf�<$t�-��������z�=�3 ��3  �   �@!�3  �-����������z���������2  ���� u�|$ u����-`��   �=�3 �G3  �   �@!�@4  Z�������̃=�P ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�Y4  ��=�P t2���\$�D$%�  =�  u�<$f�$f��f���d$u�4  ���$�2  �   ��ÍT$�=2  R��<$tmf�<$t��1  =  �?s+��������������=�3 �`2  �   �P!�]2  w:�D$��%�� D$u)��   ����-j�t�����1  ���� u�|$ u����-`��   �=�3 ��1  �   �P!��2  Z����������̃��$�1  �   ��ÍT$�h1  R��<$�D$tQf�<$t� 1  �   �u���=�3 ��1  �   �`!�1  �  �u,��� u%�|$ u����0  �"��� u�|$ u�%   �t����-`��   �=�3 �61  �   �`!�/2  Z�������U��WV�u�M�}�����;�v;���  ���   r�=�Q tWV����;�^_u�7  ��   u������r)��$���Ǻ   ��r����$��$� ��$���@d#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I ���������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���� (�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�������$�<�I �Ǻ   ��r��+��$���$�������F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I @HPX`hp��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$���������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����������������̃=�P �B8  ���\$�D$%�  =�  u�<$f�$f��f���d$�8  � �~D$f(�f(�f(�fs�4f~�fT@�f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$��4  ���D$��~D$f��f(�f��=�  |!=2  �fT ��\�f�L$�D$����f�0�fV0�fT �f�\$�D$����������������U��WV�u�M�}�����;�v;���  ���   r�=�Q tWV����;�^_u�3  ��   u������r)��$���Ǻ   ��r����$���$����$�$���#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I �tld\TLD�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�,�����$���I �Ǻ   ��r��+��$�0�$�,�@d��F#шG��������r�����$�,�I �F#шG�F���G������r�����$�,��F#шG�F�G�F���G�������V�������$�,�I ���� #�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�,��<DTh�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��;p!u���4  ��U��QQ��VW�]����  Vh?  �>  YY�M����  #�f;�uh�EQQ�$�G=  HYYtJHt9H�EWt!�`����\$�E�$jj�%<  ���HQQ�$j�;  ���7VW�I>  �E���'VW�;>  �E��E%����E��EVW�E��>  �E�YY_^������̺P��?  �P���>  ���������z�����5|>����t��j�,!  jj �xA  ���=A  jh��  j�D  Y�e� �u�N��t/��3��3�E��t9u,�H�JP����Y�v����Y�f �E������
   ��  Ë���j�mC  Y����̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�U��EV���F ��uc�G  �F�Hl��Hh�N�;8-t��*�Hpu��O  ��F;�)t�F��*�Hpu�8H  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P�Q  ��e�F�P�-P  ��Yu��P�bQ  Y��xu���M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�P  �M��E��M��H��EP�,Q  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�TB  @PV�V�������^Ë�U��j �u�d���YY]Ë�U��j �u�����YY]Ë�U���SV�u�M�������3�;�u"��  j^�0��?  �}� t�E��`p���^[��9Mv�9M~�E�3���	9Ew	�  j"��W8Mt�U3�9M��3Ƀ:-����ˋ��6����}�?-��u�-�s�} ~�N�E�����   � � F�3�8E��E��}�u����+�]h��SV��@  ����ut�N9Et�E�G�80t/�GHy���F-��d|�jd_�� F��
|�j
_�� F�� F�0@_t�90uj�APQ�q������}� t�E��`p�3������3�PPPPP�B>  ̋�U���,�p!3ŉE��ESV�uW�}j[S�M�Q�M�Q�p�0�9Q  ����u�n  ��L>  ���m�E��t���u��3Ƀ}�-��+�3Ʌ���+��M�Q�NQP3��}�-��3Ʌ�����Q�uO  ����t� ��u�E�j P�u��V�u��������M�_^3�[�����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �Y���9}}�}�u;�u#�  j^�0�i=  �}� t�E�`p����  9}v؋E��� 9Ew	�X  j"�ȋ}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW�$�������t�}� � ��  �M�ap��  �;-u�-F�} �0����$�x�Fje��V��@  YY���U  �} ���ɀ����p��@ �;  %   �3��t�-F�]������$�x����0�F�O�����  �3���'3��u$�F0�O����� ���u�U���E��  ��F1����F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~L�W#U���M�#E���� �P  f��0����9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �O  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�K�����u�E�8 u���} �4����$�p���W�@O  3�%�  #�+E�SY�x;�r	�F+����F-������ڋ��0;�|$��  ;�rSQRP�N  0�F�U�����;�u��|��drj jdRP��M  0��U�F����;�u��|��
rj j
RP��M  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u���w�ٍM�N�������u#�*  j^�0�:  �}� t�E��`p����   �} v׀} t;uu3��?-���f�0 �?-��u�-�s�G��V�^��;  @PVS�d����0�������} ~QV�^�;  @PVS�@����E����   � � ������y&�߀} u9}|�}�}������Wj0S�t������}� t�E��`p�3�_^[�Ë�U���,�p!3ŉE��EVW�}j^V�M�Q�M�Q�p�0��K  ����u�  �0��8  ���lS�]��u��  �0��8  ���S���;�t3Ƀ}�-����+��u�M�Q�M��QP3��}�-���P�J  ����t� ��u�E�j VS���N�����[�M�_3�^�/����Ë�U���,�p!3ŉE��EV�uWj_W�M�Q�M�Q�p�0�K  ����u�Q  �8�/8  ���   �M��t�S�]�3�K�}�-���<0���u��+ȍE�P�uQW�kI  ����t� �W�E�H;������|-;E}(��t
�G��u��G��u�E�j�u���u��������u�E�jP�u���u�u������[�M�_3�^�B����Ë�U��E��et_��EtZ��fu�u �u�u�u�u�'�����]Ã�at��At�u �u�u�u�u�u������0�u �u�u�u�u�u�o�����u �u�u�u�u�u�o�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3����!�����!����(r�_^Ë�Vh   h   3�V�K  ����t
VVVVV�?6  ^�j
����Q3��j ���� �� ��V�5�!�$�����u�5�3����V�5�!�(���^á�!���tP�5�3���Ѓ�!���!���tP�,���!��V6  jh ��  h���4��u�F\��f 3�G�~�~pƆ�   CƆK  C�Fh�%j�<7  Y�e� �vh�0��E������>   j�7  Y�}��E�Fl��u�8-�Fl�vl�@  Y�E������   �  �3�G�uj�6  Y�j��5  YË�VW���5�!��������Ћ���uNh  j��  ��YY��t:V�5�!�5�3���Ѕ�tj V�����YY� ��N���	V����Y3�W�8�_��^Ë�V��������uj�  Y��^�jh(�  �u����   �F$��tP�����Y�F,��tP����Y�F4��tP����Y�F<��tP����Y�F@��tP����Y�FD��tP����Y�FH��tP�u���Y�F\=�tP�d���Yj�5  Y�e� �~h��tW�<���u���%tW�7���Y�E������W   j�u5  Y�E�   �~l��t#W�?  Y;=8-t��`,t�? uW�@  Y�E������   V�����Y��  � �uj�E4  YËuj�94  YË�U��=�!�tK�} u'V�5�!�5$��օ�t�5�!�5�!���ЉE^j �5�!�5�3�����u�x�����!���t	j P�(�]Ë�Wh���4�����u	�����3�_�V�5@�h��W��h��W��3��h��W��3��h��W��3�փ=�3 �5(���3t�=�3 t�=�3 t��u$�$���3�,���3P�5�3��3� ���!�����   �5�3P�օ���   ��  �5�3�5����5�3��3���5�3��3���5�3��3�֣�3�2  ��tc�=�h�5�3���У�!���tDh  j�   ��YY��t0V�5�!�5�3���Ѕ�tj V����YY� ��N��3�@��i���3�^_Ë�U��VW3��u�0�����Y��u'9�3vV�D����  ;�3v��������uʋ�_^]Ë�U��VW3�j �u�u�F  ������u'9�3vV�D����  ;�3v��������uË�_^]Ë�U��VW3��u�u�KF  ��YY��u,9Et'9�3vV�D����  ;�3v��������u���_^]Ë�U��h ��4���th��P�@���t�u��]Ë�U���u�����Y�u�H��j��1  Y�j�1  YË�V�������V�  V��.  V�.  V�H  V�F  V�tF  ��^Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=�� th����H  Y��t
�u���Y����h,�h�����YY��uTVWhT%���������Y��;�s���t�Ѓ�;�r�=�Q _^th�Q�H  Y��tj jj ��Q3�]�j hP�Y  j��0  Y�e� 3�@94��   �4�E� 4�} ��   �5�Q�5��֋؉]Ѕ�th�5�Q�֋��}ԉ]܉}؃��}�;�rK����9t�;�r>�7�֋��r�������5�Q�֋��5�Q��9]�u9E�t�]܉]ЉE؋��}ԋ]���E�0��}�<�s�E� ��t�ЃE����E�@��}�D�s�E�� ��t�ЃE����E������    �} u)�4   j�
/  Y�u�����} tj��.  Y��k  Ë�U��j j�u������]�jj j ������Ë�U���  �u��  Yh�   ����̋�U���LV�E�P�\�j@j ^V����YY3�;�u����  ��   ��P�5�P;�s6���H��f�@� 
�Hf�@ 
�@!
�H3�H/�5�P��@�P���   ;�r�SWf9M��  �E�;��  ����E�þ   �E�;�|��9�P}k��Pj@j �����YY��tQ��P ��   �;�s1���H���` �`��`3 f�@� 
f�@ 

�@/ ���@΍P�;�r҃�9�P|����P3���~r�E�� ���t\���tW�M��	��tM��uP�X���t=����������4��P�E�� ��E�� �Fh�  �FP�T�����   �F�E�G�E�;�|�3ۋ���5�P����t���t�N��q�F���uj�X�
�C�������P�P������tB��t>W�X���t3%�   �>��u�N@�	��u�Nh�  �FP�T���t,�F�
�N@�����C���h����5�P�L�3�_[^�Ã������VW��P���t6��   ;�s!�p�~� tV�`����@   �N�;�r��7�����' Y�����Q|�_^Ã=�Q u�_6  V�5�3W3���u����   <=tGV�[-  Y�t���u�jGW�������YY�=�3��tˋ5�3S�3V�*-  �>=Y�Xt"jS����YY���t?VSP�,  ����uG���> u��5�3������%�3 �' ��Q   3�Y[_^��5�3������%�3 �����3�PPPPP�3*  ̋�U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�3D  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�NC  Y��t��M�E�F��M��E���+C  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9�Qu��3  h  �4VS�5�d���Q�5�3;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�������Y;�t)�U��E�P�WV�}�������E���H��3�5�33�����_^[�Ë�U���SV�p���3�;�u3��wf93t��f90u���f90u�W�=l�VVV+�V��@PSVV�E��׉E�;�t8P�;���Y�E�;�t*VV�u�P�u�SVV�ׅ�u�u������Y�u�S�h��E��	S�h�3�_^[�Ë�V�p�pW��;�s���t�Ѓ�;�r�_^Ë�V�x�xW��;�s���t�Ѓ�;�r�_^�j h   j �t�3Ʌ����5����55�x��%5 �����h&d�5    �D$�l$�l$+�SVW�p!1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35p!W��E� �E�   �{���t�N�38�8����N�F�38�(����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t����)  �E���x@G�E��؃��u΀}� t$����t�N�38�����N�V�3:�����E�_^[��]��E�    �ɋM�9csm�u)�=�P t h�P�>  ����t�UjR��P���M�U�t)  �E9Xthp!W�Ӌ��v)  �E�M��H����t�N�38�����N�V�3:�����E��H���
)  �����9S�O���hp!W���!)  ������U��V����������2  �N\�U��W9t�����   ;�r���   ;�s9t3���t�P��u3���   ��u�` 3�@��   ����   �MS�^`�N`�H����   j$Y�~\�d9 �����   |� �~d=�  �u	�Fd�   �~=�  �u	�Fd�   �n=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=� �u	�Fd�   �=� �u�Fd�   �vdj��Y�~d��` Q��Y�^`[���_^]Ë�U��csm�9Eu�uP����YY]�3�]Ë�U����p!�e� �e� SW�N�@��  ��;�t��t	�Уt!�eV�E�P����u�3u����3�� �3����3��E�P�|��E�3E�3�;�u�O�@����u��G  ����5p!�։5t!^_[�Ë�U��} u�-  �    �#  ���]��uj �55���]�f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U�����U��3��M;�8�t
@��r�3�]Ë�<�]Ë�U����  �p!3ŉE�SV�uWV������3�Y�����;��l  j�!?  Y���  j�?  Y��u�=�3��   ���   �6  ht�h  � 5W�z>  ������   h  �R5VSf�Z7�����  ��uhD�SV�B>  ����t3�PPPPP��   V�>  @Y��<v*V�>  �E�4��+�j��h<�+�SP�=  ����u�h4��  VW�<  ����u������VW�v<  ����u�h  h��W��:  ���^SSSSS�y���j��P���;�tF���tA3��G�����f9Gt@=�  r�S�����P�����P�]��"  YP�����PV����M�_^3�[������j�=  Y��tj�=  Y��u�=�3uh�   �%���h�   ����YYË�U��E3�;��!tA��-r�H��wjX]Ë��!]�D���jY;��#���]�������u�X#Ã��������u�\#Ã�Ë�U��V������MQ�����Y�������0^]Ë�U��E�H;]Ë�U���5H;����t�u��Y��t3�@]�3�]�j
����P3�����������������U�������$�~$�   ��fD$f��f%�f-00f=��B  f���Y�f���-��X�f��\�f( ��Y�fɁ�v ����?f(-��������fY��\��Y��\�fxf����\�fY�f\�f(5���Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-���Y fX5��fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f@��\�fL$�D$��������I ���̀zuf��\���������?�f�?f��^���٭^����|��剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����|��剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����t����۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-`���p��� ƅp���
��
�t�����������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   ��   Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t�{   Z��]   Z��,$Z����������������������   s��������������������������   v���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�7  ���E�f�}t�m���������������U�������$�~$�   ��fD$f%��f��fW�f����fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU��fV�f($������X��\��Y��Y��Y����X��^�f=8�f-(��\�fs�?��fs�?�Y�fp�Df50��Y��Y���fW��Y��Y��X��Y��X�fp���X��X��X�fD$�D$���-�  ��C�  �Y��\��Q�f��fs�fT= �fs���f%�����\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<����Y�f(���Y��Y��\��X��\��X�f-(��\��X�f8��^�f0�f\������Y�%�   ���Y��Y΃��Y��Y��X�f���Y��X�f���X�fp���\��X�fV�fD$�D$����;  = 8  sjf�f(5@�f�f(P�f(%`�fY���fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X�fD$�D$���-�;  ���O  �Y��\��Q�f��fT=�fp�DfT���f%�����\��Y��X��Y��\����Y��Y��\��\��X��\�f(@�fp���\��X�fp���X��Y��X�fp���^�f(p�f(-P�f(`�fY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f(���Y�fX�fp���Y��fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fV�fD$�D$����� = � ��   f~�fs� f~�����  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$�  fD$����fD$�D$���f��f��f���X�fU�fV���fD$�D$���fD$fW��Xƺ�  �t���fD$fW�����f�����  �����  r�X�fV��Y�fD$�D$���W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y������U���(3��E��E�9P;t�5�P�����k�M��   V;���  ��  ���  �  jZ+���   I��   ����   I��   ����   ItN��	�  �E�   �E�|��M��M�u�]���M��]�Q��]���Y����  ����� "   ��  �E�x��M��M�u�]���M��]�Q��E�   �]���Y�  �E�   �E�x���E�p��M�u��M�]���]���?  �U��E�p��W����E�l��ΉU��E�l��?����E�|��q�����tWItHIt9It ��t���  �E�d���E�\���E�|��M��u��u����E�|��c����E�   �������E���   �E�   �E�T��������������   �$�<�E�l���E�p���E�x���E�L���E�D��t����E�<��h����E�4��\����E�0���E�,���E�(��M��u�M����M�]���]�M��]�Q�E�   ��Y��u������ !   �E��^�Ðg;p;y;�;�;�;;�;�:�:�;�;�;��U��QQSV���  V�5`#�  �EYY�M�ظ�  #�QQ�$f;�uU�	  YY��~-��~��u#�ESQQ�$j�0  ���tVS�
  �EYY�f�ES�`����\$�E�$jj�A��.  �]��E�Y�EY������DzVS�v
  �E�YY�"�� u��E�S���\$�E�$jj�  ��^[�Ë�U���(  �`<�\<�X<�T<�5P<�=L<f�x<f�l<f�H<f�D<f�%@<f�-<<��p<�E �d<�E�h<�E�t<��������;  �h<�d;�X;	 ��\;   �p!�������t!�����������;j��-  Yj ���h������=�; uj�-  Yh	 ����P����Ë�U��� �e� Wj3�Y�}��9Eu�����    �}  ����x�MV�u��t��u�����    �Y  ����S�����E�;�w�M��u�E��u�E�B   �u�u�P�u��/  ������t�M�x�E��  ��E�Pj ��,  YY��^_�Ë�U���uj �u�u�u�<�����]Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u����M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�  Y����  �t�Etj�e  Y����x  ����   �E��   j�C  �EY�   #�tT=   t7=   t;�ub��M����`$��{L�H��M�����{,�`$�2��M�����z�`$���M�����z�P$��P$��������   ���   �E��   3��t��W�}���������D��   ��E�PQQ�$�l  �M��]�� �����������}�E���H��S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}� ���� "   ]������� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���h#;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�'  ����uV�,���Y�E�^�Ë�l#�h��  �u(�  �u�����E ���Ë�U��=@- u(�u�E���\$���\$�E�$�uj�/�����$]������h��  �u� !   �H  �EYY]Ë�S��QQ�����U�k�l$���   �p!3ŉE��s �CP�s��������u#�e��P�CP�CP�s�C �sP�E�P�j������s�o������=@- u+��t'�s �C���\$���\$�C�$�sP�q�����$�P�����$��  �s �  �CYY�M�3�������]��[Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]�f�M��  V��f#�^f;�uj���  f;�u�E�� u9Utj��3�]Ë�U���E������������Dz3��   �E3ɩ�  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������&Q���EQQ�$������U�����  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��f#E�f����E�m�E��Ë�U��QQ�M��t
�-x$�]���t����-x$�]�������t
�-�$�]����t	�������؛�� t���]����jhp�����3�9�QtV�E@tH9�$t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�$ �e��U�E�������e��U����������������U���0���S�ٽ\�����=@- t������8����   [����ݕz������U���U���0���S�ٽ\����=@- t�s�����8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8��������   [�À�8�����=�3 uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ������������������s4�(��,ǅr���   ������������� �����v� �VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P��  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8������������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[���  ��tj�  Y��$tjh  @j�J   ��j����̋�U��M��$�U#U��#�ʉ�$]Ë�U��E�|>]Ë�U��E��>]Ë�U���(  �p!3ŉE�S�]W���tS�8   Y������ jL������j P�h�����������������0�����������������������������������������������f������f������f������f������f������f��������������E�M������ǅ0���  �������I��������M�������M���������������j �����������P�����u��u���tS�C  Y�M�_3�[�����Ë�Vj� �Vj�������V���P���^Ë�U���5�>����t]���u�u�u�u�u�����3�PPPPP�������Ë�VW3���>�<��$u���$�8h�  �0���T���tF��$|�3�@_^Ã$��$ 3����S�`�V��$W�>��t�~tW��W蹯���& Y�����%|ܾ�$_���t	�~uP�Ӄ����%|�^[Ë�U��E�4Ũ$���]�jh�����3�G�}�3�95u����j����h�   �s���YY�u�4��$9t���mj�N���Y��;�u������    3��Pj
�X   Y�]�9u+h�  W�T���uW����Y������    �]���>�W�ͮ��Y�E������	   �E������j
�)���YË�U��EV�4Ũ$�> uP�#���Y��uj�9���Y�6���^]Ë�U��UVW��t�}��u�D���j^�0�������3�E��u����+���@��tOu��u� ����j"Y�����3�_^]��������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�������SVW�T$�D$�L$URPQQhPd�5    �p!3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�R+  �   �C�d+  �d�    ��_^[ËL$�A   �   t3�D$�H3��Q���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�*  3�3�3�3�3���U��SVWj Rh�PQ�<l  _^[]�U�l$RQ�t$������]� ��������������U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP蝪��3��ȋ��~�~�~����~�����%���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �p!3ŉE�SW������P�v����   ����   3�������@;�r�����ƅ���� ��t0���������;�w+�@P������j R�ک�����C����u�j �v�������vPW������Pjj �8,  3�S�v������WPW������PW�vS��*  ��DS�v������WPW������Ph   �vS��*  ��$3���E������t�L���������t�L ��������  ���  @;�r��R��  ǅ��������3�)�������������  ЍZ ��w
�L�Q ���w�L �Q����  A;�rƋM�_3�[�S�����jh��t�����������*�Gpt�l t�wh��uj �O���Y�������j�����Y�e� �wh�u�;5�)t6��tV�<���u���%tV�]���Y��)�Gh�5�)�u�V�0��E������   뎋u�j����YË�U���S3�S�M�谶���@���u�@   ���8]�tE�M��ap��<���u�@   ����ۃ��u�E��@�@   ��8]�t�E��`p���[�Ë�U��� �p!3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9� *��   �E��0=�   r����  �t  ����  �h  ��P������V  �E�PW������7  h  �CVP�����3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP趦���M��k�0�u���*�u��+�F��t)�>����E����)D;�FG;�v�}���> uЋu��E����}��u�r�ǉ{�C   �i���j�C�C��*Zf�1f�0����Ju������������L@;�v����~� �0����C��   �@Iu��C�����C�S��s3��ȋ�����{����95@�T�������M�_^3�[�J�����jh��k����M���������}�������_h�u�q����E;C�W  h   ����Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�<���u�Fh=�%tP�5���Y�^hS�=0����Fp��   ��*��   j�\���Y�e� �C�$@�C�(@�C�,@3��E��}f�LCf�E@@��3��E�=  }�L���'@��3��E�=   }��  ���(@���5�)�<���u��)=�%tP�|���Y��)S���E������   �0j�����Y��%���u ���%tS�F���Y�#����    ��e� �E��#���Ã=�Q uj��V���Y��Q   3�Ë�U��SV�50�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��*t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5<�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��*t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�U��SV�u���   3�W;�to=h-th���   ;�t^9uZ���   ;�t9uP襣�����   �7)  YY���   ;�t9uP脣�����   �(  YY���   �l������   �a���YY���   ;�tD9u@���   -�   P�@������   ��   +�P�-������   +�P�������   ���������   =�*t9��   uP�$  ���   ����YY�~P�E   ���*t�;�t9uP�Ƣ��Y9_�t�G;�t9uP询��Y���Mu�V蠢��Y_^[]Ë�U��W�}��t;�E��t4V�0;�t(W�8�j���Y��tV������> Yu��`,tV�s���Y��^�3�_]�jh�������5������*�Fpt"�~l t�����pl��uj �����Y�������j�Y���Y�e� �58-��lV�Y���YY�E��E������   �j�R���Y�u�Ë�U����u�M��[����E����   ~�E�Pj�u�B(  ������   �M�H���}� t�M��ap��Ë�U��=l@ u�E�(-�A��]�j �u����YY]Ë�U���SV�u�M��ڮ���]�   ;�sT�M胹�   ~�E�PjS�'  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�(  YY��t�Ej�E��]��E� Y������ *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�   ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=l@ u�E�H���w�� ]�j �u�����YY]Ë�U���(�p!3ŉE�SV�uW�u�}�M�舭���E�P3�SSSSW�E�P�E�P�2  �E�E�VP�g'  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�����Ë�U���(�p!3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P�n1  �E�E�VP�,  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�I����Ë�U��MS�YV�u3�;�u����j^�0�g������   9Ev�U�;�~��@9Ew�`���j"Y�����W�~�0�ǅ�~���t��C�j0Y�@J���M�  ��x�;5|�� 0H�89t�� �>1u�A�W����@PWV蝡����3�_^[]Ë�U��Q�M�AS����% �  V��  #�W�E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��B��<  �U����������U��E����������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0�p!3ŉE��ES�]V�E�W�EP�E�P�"���YY�E�Pj j���uЋ���f��46  �u܉C�E��E��C�E�P�uV�}�����$��u�M�_�s^��3�[�b�����3�PPPPP�G������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�z���YË�U��E�M%����#�V�u������t$��tj j ��>  YY��u���j^�0�P������P�u��t	�>  ���>  YY3�^]Ë�U��M��tj�3�X��;Es�-����    3�]��MV���uF3����wVj�55����u2�=L; tV�F���Y��uҋE��t�    3���M��t�   ^]Ë�U��} u�u�>���Y]�V�u��u�u迚��Y3��MW�0��uFV�uj �55�������u^9L;t@V�����Y��t���v�V����Y�Y����    3�_^]��H�������P�����Y����0�������P�����Y�����jh������ ����@x��t�e� ���3�@Ëe��E����������������h�b���4@Ë�U��E�8@�<@�@@�D@]Ë�U��E���V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5@@���j h0�2���3��}�}؋]��Kt��jY+�t"+�t+�tY+�uC�Գ�����}؅�u����T  �8@�8@�U�w\���]���Y�p��Q�Ã�t2��t!Ht������    �����빾@@�@@��<@�<@�
�D@�D@�E�   P���E�3��}���   9E�uj�F���9E�tP� ���Y3��E���t
��t��u�O`�MԉG`��u>�Od�M��Gd�   ��u,����M܋����9M�}�M�k��W\�D�E���葱����E������   ��u�wdS�U�Y��]�}؃}� tj ����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3������Ë�U��E�L@]������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��t�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�hPh&d�    P��SVW�p!1E�3�P�E�d�    �e��E�    h   �*�������tT�E-   Ph   �P�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE�3ҁ9  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U����u�M��	����E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U���$�p!3ŉE��ES�E��EVW�E��:����e� �=P@ �E�u}h����؅��  �=@�hS�ׅ���   �5�P��h�S�P@��P��h�S�T@��P��h�S�X@��P�֣`@��th�S��P�֣\@�\@�M�5�;�tG9`@t?P���5`@���֋؅�t,��t(�ׅ�t�M�Qj�M�QjP�Ӆ�t�E�u	�M    �3�T@;E�t)P�օ�t"�ЉE��t�X@;E�tP�օ�t�u��ЉE��5P@�օ�t�u�u��u��u����3��M�_^3�[�0����Ë�U��V�uW��t�}��u�t���j^�0�O�����_^]ËM��u3�f��݋�f�: t��Ou��t�+��f�
��f��tOu�3���u�f��"���j"Y���몋�U��US�]VW��u��u9Uu3�_^[]Å�t�}��u�����j^�0��������݅�u3�f��ЋM��u3�f��ԋ��u��+��f���f��t'Ou��"��+��f���f��tOtKu��u3�f����y���3����u�MjPf�DJ�X�d���f��X���j"Y����j�����U��Ef���f��u�+E��H]Ë�U��V�uW��t�}��u����j^�0�������_^]ËE��uf��ߋ�+��f���f��tOu�3���u�f������j"Y���뼋�U��M��x��~��u��3]á�3��3]������    �y������]Ë�S��QQ�����U�k�l$���   �p!3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|������������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�z�����h��  ��x��������>YYt�=@- uV�    Y��u�6�L���Y�M�_3�^�������]��[�3�Ë�U��QQ�E���]��E��Ã%�P Ë�U��QV�uV�&C  �E�FY��u����� 	   �N ����/  �@t������ "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�A  �� ;�t��@  ��@;�u�u�@  Y��uV�>@  Y�F  W��   �F�>�H��N+�I�N;�~WP�u�:?  ���E��M�� �F����y�M���t���t������������P���!�@ tjSSQ�7  #����t%�F�M��3�GW�EP�u��>  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��QSV����艿���G@� �E�t
� u�J�o����  �(�E� ��K�����E�>�u�P����8*u�ϰ?�u�������9����8 u
�/����M��^[�Ë�U���x  �p!3ŉE�S�]V�u3�W�u�}�������������������������������������������������������������v�����u+趾���    ���������� t
�������`p������
  �F@u^V�@  Y��!���t���t�ȃ���������P����A$u����t���t�ȃ�������P����@$��q���3�;��g����3ɉ��������������������������9
  G������9������&
  �B�<Xw���� ���3����@j��Y������;���	  �$�Gy��������������������������������������������	  �� tJ��t6��t%HHt���u	  �������i	  �������]	  �������Q	  �������   �B	  �������6	  ��*u,���������[�������;��	  �������������	  ������k�
�ʍDЉ�������  ��������  ��*u&���������[�������;���  ��������  ������k�
�ʍDЉ������  ��ItU��htD��lt��w��  ������   �r  �?luG������   �������W  �������K  ������ �?  �<6u�4u�������� �  �������  <3u�2u�������������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������ ������P��P�  Y��������Yt"�����������������G������������������������������h  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@�������   ������������9������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  �������[���������  ;�u�H-������������ǅ����   �y  ��X��  HHty+��'���HH��  ��������  ������t0�C�Ph   ������P������P�=  ����tǅ����   ��C�������ǅ����   �������������/  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  �D-������P�u���Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�3���������(;  ���:��������� tf������f���������ǅ����   ��  ������@ǅ����
   �������� �  ��  ��S����  u��gucǅ����   �W9�����~�������������   ~=��������]  V袦��������Y��������t���������������
ǅ�����   ��5����������C�������������P��������������������P������������WP�5�!���Ћ���������   t������ u������PW�5�!����YY������gu��u������PW�5�!����YY�?-u������   G������W�
���ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �p���������Qƅ����0������ǅ����   �L�����   �R������� t��������@t�C���C����C���@t��3҉�������@t��|��s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW��  ��0���������ڃ�9~������N뽍E�+�F������   ������������tb��t�΀90tW�������������0@�?If90t��;�u�+��������(;�u�D-�������������I�8 t@;�u�+����������������� �}  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+������������u'����~!������������� O�F����������t��ߋ�����������������P�������N���������Yt(������u��������ϰ0K������������t��ヽ���� ������tT��~P�������Pj�E�P������PK���8  ����u ��������t�E�P�����������Y��u����������������������������Y������ |.������t%��������������ϰ K�H����������t��ヽ���� t���������������� Y���������������t������������3�������������� t
�������`p��������M�_^3�[�?����ÍI 2q1oao�opp\p�q��U��E��t���8��  uP�z���Y]����������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� �����������U��SVWUj j hHz�u�B  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�hPzd�5    �p!3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �yPzu�Q�R9Qu�   �SQ�P-�SQ�P-�L$�K�C�kUQPXY]Y[� ��Ë�U����p!3ŉE��US3�VW;�~�E��I8t@;�u������+�H;�}@�E�]�9]$u�E� �@�E$�5��3�9](SS�u���u��   P�u$�֋��}�;�u3��R  ~Cj�3�X����r7�D?=   w�4  ��;�t� ��  �P�N���Y;�t	� ��  ���E���]�9]�t�W�u��u�uj�u$�օ���   �5��SSW�u��u�u�։E�;���   �   �Mt)�E ;���   9E���   P�uW�u��u�u���   �}�;�~Bj�3�X����r6�D?;�w��3  ��;�th���  ���P���Y;�t	� ��  �����3�;�t?�u�W�u��u��u�u�օ�t"SS9] uSS��u �u�u�WS�u$�l��E�W�8���Y�u��/����E�Y�e�_^[�M�3��5����Ë�U����u�M��7����u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap��Ë�U��QQ�p!3ŉE�S3�VW�]�9]u�E� �@�E�5��3�9] SS�u���u��   P�u�֋�;�u3��~<�����w4�D?=   w�2  ��;�t� ��  �P�R~��Y;�t	� ��  ���؅�t��?Pj S�}����WS�u�uj�u�օ�t�uPS�u����E�S�����E�Y�e�_^[�M�3������Ë�U����u�M��
����u$�E��u�u�u�u�uP��������}� t�M��ap��Ë�U��V�u���c  �v�*~���v�"~���v�~���v�~���v�
~���v�~���6��}���v ��}���v$��}���v(��}���v,��}���v0��}���v4��}���v��}���v8�}���v<�}����@�v@�}���vD�}���vH�}���vL�}���vP�}���vT�}���vX�x}���v\�p}���v`�h}���vd�`}���vh�X}���vl�P}���vp�H}���vt�@}���vx�8}���v|�0}����@���   �"}�����   �}�����   �}�����   �}�����   ��|�����   ��|�����   ��|�����   ��|�����   ��|�����   �|�����   �|�����   �|�����   �|�����   �|�����   �|�����   �}|����@���   �o|�����   �d|�����   �Y|�����   �N|�����   �C|�����   �8|�����   �-|�����   �"|�����   �|�����   �|�����   �|�����   ��{�����   ��{����   ��{����  ��{����  ��{����@��  �{����  �{����  �{����  �{����  �{����   �{����$  �z{����(  �o{����,  �d{����0  �Y{����4  �N{����8  �C{����<  �8{����@  �-{����D  �"{����H  �{����@��L  �	{����P  ��z����T  ��z����X  ��z����\  ��z����`  ��z����^]Ë�U��V�u��tY�;h-tP�z��Y�F;l-tP�z��Y�F;p-tP�z��Y�F0;�-tP�yz��Y�v4;5�-tV�gz��Y^]Ë�U��V�u����   �F;t-tP�Az��Y�F;x-tP�/z��Y�F;|-tP�z��Y�F;�-tP�z��Y�F;�-tP��y��Y�F ;�-tP��y��Y�F$;�-tP��y��Y�F8;�-tP��y��Y�F<;�-tP�y��Y�F@;�-tP�y��Y�FD;�-tP�y��Y�FH;�-tP�{y��Y�vL;5�-tV�iy��Y^]Ë�U���S�u�M������]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�X����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M��4����E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���8�p!3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=�-O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC��-��+�-;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5�-N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3���-�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  ��-;�-��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy��-�-3�@�   �-�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+�-��M���Ɂ�   �ً�-]���@u�M̋U�Y��
�� u�M̉�M�_3�[�~���Ë�U���8�p!3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=�-O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC��-��+�-;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5�-N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3���-�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  ��-;�-��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy��-�-3�@�   �-�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+�-��M���Ɂ�   �ً�-]���@u�M̋U�Y��
�� u�M̉�M�_3�[�Ey���Ë�U���|�p!3ŉE��E3�V3��E��EFW�E��}��M��u��M��M��M��M��M��M��M�9M$u�V����    �0���3��<  �U�U��< t<	t<
t<uB��S�0�B���  �$���Hπ�wjYJ�ߋM$�	���   �	:ujY������+tHHt���|  ���jY�E� �  뤃e� jY뛍Hωu���v��M$�	���   �	:uj�<+t"<-t:�t�<C�/  <E~
,d<�!  j�Jj넍Hπ��_����M$�	���   �	:�a���:��s����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�h���<+t�<-t��k����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Hπ�wj	��������+t HHt���=���j�����M��jY�Q���j�~����u���B:�t�,1<v�J�&�Hπ�v�:�뿃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�]����B:�}��Q����M��E�O�? t�E�P�u��E�P�  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �!  =�����-  ��0��`�E�;���  }�ع�1�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k��� �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��   f;��  ���  f;��	  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� ����E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��yB��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  f9E�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �=����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W[�M�_3�^�r���ÍI Ώ �k�����-���q�������U���t�p!3ŉE��E�U� �  #�S�]�E��A�V#�f�}� W�]��E������E������E����?�E�   t�C-��C �u�}f��u7����   ����   3�f9M�f�����$ �Cf�C0�C 3�@�  f;���   �M3�@f��   �;�u�} t��   @uh@�S3�PPPPP�}���3�f9U�t��   �u9Uu-h8�;�u"9Uuh0�CjP�W�������u��C�h(�CjP�:�������u��C3��k  �ʋ�i�M  �������Ck�M��������3�f�M��ع�0��`�ۉE�f�U�u�}�M���  ��y��1��`�ۉE�����  �E�T�������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E����E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��yB��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��}����M�����?  ��  f;���  �]��E�3҉U��U��U�U��U�3�#�#Ё� �  �4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��Z���3�3�f9u���H%   � ���E��a���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~K�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m����M��}� ����E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��yB��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t0����)3�f�� �  f9E�f�B0����$ �B�B �s�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�y2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K����C���<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[�i���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}�f�]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   �é   t��   �}�M����#�#���E;���   ���������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95�Q��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��M���Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[�Ë�U��QQ�EV�u�E��EWV�E��Z  ���Y;�u�d���� 	   �ǋ��J�u�M�Q�u�P����E�;�u����t	P�V���Y�ϋ������P�����D0� ��E��U�_^��jhp�́������]܉]��E���u������  ������ 	   �Ë��   ��x;�Pr�ӈ���  踈��� 	   蒨���ы����<��P��������L1��t�P��  Y�e� ��D0t�u�u�u�u��������E܉U���V���� 	   �^����  �]܉]��E������   �E܋U��?�����u�  YË�U���  �  �p!3ŉE��EV�uW3���4�����8�����0���9}u3��  ;�u�����8�χ���    詧������  ������S���P������L8$�����$�����?�����t��u'�M����u苇���  �p����    �J����  �D8 tjj j V������V�>  Y����  ��D���  �?r���@l3�9H�� �����P��4�����3�;��`  ;�t8�?����P  �����4����� ���3���,���9E�#  ��@�����?������g  ���$���3���
��������ǃx8 t�P4�U�M��`8 j�E�P�K��P�#���Y��t:��4���+�M3�@;���  j��D���SP��  �������  C��@����jS��D���P�  ������n  3�PPj�M�Qj��D���QP�� ���C��@����l������=  j ��,���PV�E�P��$���� �4������
  ��@�����0������8���9�,�����  ����� ��   j ��,���Pj�E�P��$���� �E��4�������  ��,�����  ��0�����8����   <t<u!�33Ƀ�
������@�����D��������<t<uR��D����.  Yf;�D����I  ��8�������� t)jXP��D����  Yf;�D����  ��8�����0����E9�@���������  ����8����T4��D8��  3ɋ�D8���  ��?��� ��D�����   ��4���9M��  ��3�+�4�����H���;Ms&�CA�� �����
u��0���� @F�@F���  rՋ���H���+�j ��(���PV��H���P��$���� �4������C  ��(����8���;��;  ��+�4���;E�l����%  ��?�����   ��4���9M�H  ��@��� ��+�4���j��H���^;MsC��Ή� �����
u�0���j[f��� �����@����@���f�Ɓ�@����  r�����H���+�j ��(���PV��H���P��$���� �4������i  ��(����8���;��a  ��+�4���;E�G����K  ��4�����,���9M�u  ��,�����@��� +�4���j��H���^;Ms;��,�����,���΃�
uj[f���@����@���f�Ɓ�@����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �l���;���   j ��(���P��+�P��5����P��$���� �4�����t�(���;�������D���;�\��,���+�4�����8���;E�����?Q��(���Q�u��4����48�����t��(�����D��� ��8��������D�����8��� ul��D��� t-j^9�D���u葁��� 	   虁���0�?��D���蝁��Y�1��$���� �D@t��4����8u3��$�Q����    �Y����  ������8���+�0���[�M�_3�^��\����jh���y���]���u�����  ����� 	   ����   ��x;�Pr������  �ۀ��� 	   赠���ҋ����<��P�������D0��t�S��  Y�e� ��D0t�u�uS�n������E��聀��� 	   艀���  �M���E������   �E��oy��Ë]S�B  YË�U���p@h   �n��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u����� 	   3�]Å�x;�Pr����� 	   賟���ދȃ������P���D��@]ø�-á�PVj^��u�   �;�}�ƣ�PjP�n��YY��@��ujV�5�P��m��YY��@��ujX^�3ҹ�-���@��� ����x0|�j�^3ҹ.W�������P����������t;�t��u�1�� B��h.|�_3�^���
  �= 4 t�  �5�@��N��YË�U��V�u��-;�r"��X0w��+�����Q�����N �  Y�
�� V���^]Ë�U��E��}��P�����E�H �  Y]ËE�� P���]Ë�U��E��-;�r=X0w�`���+�����P�Ϟ��Y]Ã� P���]Ë�U��M�E��}�`�����Q蠞��Y]Ã� P���]Ë�U��E��u��}���    �ĝ�����]Ë@]áp!��3�9t@����Ë�U���SV�u3�W�};�u;�v�E;�t�3��{�E;�t�������v�}��j^�0�[������V�u�M��[���E�9X��   f�E��   f;�v6;�t;�vWSV�LL�����5}��� *   �*}��� 8]�t�M��ap�_^[��;�t&;�w �
}��j"^�0����8]�t��E��`p��y�����E;�t�    8]��<����E��`p��0����MQSWVj�MQS�]�p�l�;�t9]�j����M;�t�������z�P���;��s���;��k���WSV�K�����[�����U��j �u�u�u�u������]�������������Q�L$+ȃ����Y�  Q�L$+ȃ����Y�  ����U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U����ES3�VW�E�N@  ��X�X9]�E  �]����}襥��э<	���ʋU�e ��ى}����֋u����ϋ��M���U�����։0�x�H;�r;U�s�E   �} �t'�u��e �~;�r��s�E   �} �xtA�H�u�e �7;�r;�s�E   �} �XtA�HM��e� ��ɋ��������މH�M�M�M��X�1�2�u�;�r;�s�E�   �}� �t$�K3�;�r��s3�B�ىH��t
�M�A�M�H�M�M�E�} �X�H�����3�9Xu*�P��E���  ��������������P�;�t܉x�x�� �  u0�H��E���  �����������ʉ�H�x�� �  t�f�M�_^f�H
[�Ë�U��MS3�VW;�|[;�PsS��������<��P����D0t6�<0�t0�=�3u+�tItIuSj��Sj��Sj�������3���,y��� 	   �4y������_^[]Ë�U��E���u�y���  ��x��� 	   ���]Å�x;�Pr��x���  ��x��� 	   賘���Ջ������P�����Dt͋]�jh��qq���}����������4��P�E�   3�9^u5j
����Y�]�9^uh�  �FP�T���u�]��F�E������0   9]�t�����������P�D8P����E��2q���3ۋ}j
觘��YË�U��E�ȃ������P���DP���]Ë�U��Q�=P3�u��  �P3���u���  ��j �M�Qj�MQP�����t�f�E�Ë�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��$U���E�9Xu�E;�t�f�8]�t�E��`p�3�@�ˍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p������E�u�M;��   r 8^t���   8]��f����M��ap��Z�����v��� *   8]�t�E��`p�����;���3�9]��P�u�E�jVj	�p������:���뺋�U��j �u�u�u�������]������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��jh��	o��3ۉ]�j蝗��Y�]�j_�}�;=�P}T����@9�tE���@�tP��  Y���t�E��|(��@���� P�`���@�4���E��Y��@��G��E������	   �E���n���j�B���YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�{���YP�L�����;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV����P�A  Y��Y��3�^]�jh��m��3��}�}�j�N���Y�}�3��u�;5�P��   ��@��98t^� �@�tVPV����YY3�B�U���@���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��uࡀ@�4�V� ���YY��E������   �}�E�t�E��>m���j踔��Y�j����Y������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� 3�PPjPjh   @hH����P3áP3���t���tP���Ë�U��V�uW�����u�s���    �k�����D�F�t8V�����V���N  V�m���P�~  ����y�����F��tP�fC���f Y�f ��_^]�jh��k���M��3��u������u�s���    ���������F@t�f �E��	l���V����Y�e� V�<���Y�E��E������   �ԋuV�b���Y�jh8�k���]���u�r��� 	   ����   ��x;�Pr�r��� 	   �h����ڋ����<��P�������D��t�S����Y�e� ��Dt1S�0���YP�����u���E���e� �}� t�4r���M��r��� 	   �M���E������   �E��k��Ë]S�����Y�������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U��V�uWV�Y���Y���tP��P��u	���   u��u�@Dtj�.���j���%���YY;�tV����YP�����u
�����3�V�u����������P����Y�D0 ��tW�q��Y����3�_^]�jhX�i���]���u��p���  ��p��� 	   ����   ��x;�Pr�p���  �p��� 	   �v����ҋ����<��P�������D0��t�S����Y�e� ��D0tS�����Y�E���Jp��� 	   �M���E������   �E��@i��Ë]S����YË�U��V�u�F��t�t�v�!@���f����3�Y��F�F^]��%����������U��`3�a��h@��>����]�����U��j �|3豨��]����������������U��`3�a��]�                                                                                                                                                                                 � � � � � �   , 8 F T ^ v � � � � � � � � $ 2 D \ r � � � � � �   2 > J ` t � � � � �    $ 0 : F X f v � � � � � � �             � �        ^�7a-�W7�        #��                    �������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?Ocontainer.png  Ocontainer      �  � @ p � @ � 0; P; `; @; �; �; �; �; p; �; �M �M O `O �P �Q  R �Q �Q �Q �Q �Q �Q PO 0O @O              �o@333333�?      �?ffffff�?src/ContainerObject.cpp ../../resource/_api/c4d_resource.cpp    #   #   #   #   #   #   #   #   #   #   M_EDITOR    M_EDITOR    �P: �������N���������������C-DT�!	@-DT�!�?res     �������N���������������C-DT�!	@-DT�!�?�������?-DT�!��      �-DT�!�?      Y@�������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_misc/datastructures/basearray.h      �������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ~   Progress Thread 0%  ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp %   ../../resource/_api/c4d_gui.cpp �� � � � 0� @� P�  � 0�     �������������     �f@-DT�!	@     @�@X� � � � 0� @� P�  � P� �p� `� p� �  � �� �� 0� �� @�  � � � � � � 0� @� P�  �  � 8p� � � � 0� @� P�  � �� �� ��  � �  � 0� @� P� �� � �� �� �������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_file.cpp    ../../resource/_api/c4d_file.cpp    �������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ����MbP?��I�8   %s      c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_general.h    �������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp          �?  4&�k�  4&�kC �Ngm��C   ����A�`�P�r	r	../../resource/_api/c4d_pmain.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ��`�              �?      �?3      3            �      0C       �       ��              fmod         d	�0o0�040�0o0�0m0m0�0m0�0�0o0�0e+000   K E R N E L 3 2 . D L L     FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �      r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            ��   ��	   (�
   ��   ��   (�   ��   ��   �   ��   X�   ��   ��   X�   ��    (�!   8�x   �y   ��z   ���   ���   ��M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y     
 
     . . .   < p r o g r a m   n a m e   u n k n o w n >     R u n t i m e   E r r o r ! 
 
 P r o g r a m :                                           �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������               ���5�h!����?      �?            �?5�h!���>@�������             ��      �@      �                          8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �              �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow X;�;_nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    �������             ��      �@      �         Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        ��������������|�t�h�\�Y�T�L�H�D�@�<�8�4�0�$� �������� ���������������������������������������������������|�d�X�D�$����������d�@� �����������������x�h�L�,��������l�H�$�������Y�����l�L�0�H H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L     ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx                                                                                                                                                                                                                                                                                                ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ 1#QNAN  1#INF   1#IND   1#SNAN  C O N O U T $   ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           p!`              8             ����    @             ����    @   T           d8               |�8    0        ����    @   l            L �           ���8    L        ����    @   �             T            l $           4<    l         ����    @   $            � l           |�<    �        ����    @   l            � �           ��    �         ����    @   �            �             <    �        ����    @                � L           \l<    �        ����    @   L            � �           ��    �         ����    @   �            !�           ��    !        ����    @   �             !,           <D     !        ����    @   ,& P Pz                     ����    ����    ����    �    ����    ����    ����b�s�    ����    ����    ����    ��    ����    ����    ����    
    ����    ����    ����    f����    u����    ����    ����    (����    4����    ����    ����    v    ����    ����    ����H,H    ����    ����    ����    GN    ����    ����    ����    �S    ����    ����    ����    �W    ����    ����    ����    [    ����    ����    �����b�b    ����    ����    ����    �d    ����    ����    ����Kf^f    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    Ĵ    ����    ����    ����    .�    ����    ����    ����    ��        ������    ����    ����    �    ����    ����    ����    �    ����    ����    ����    ���         2  �                     � � � � � �   , 8 F T ^ v � � � � � � � � $ 2 D \ r � � � � � �   2 > J ` t � � � � �    $ 0 : F X f v � � � � � � �        �GetCurrentThreadId  � DecodePointer �GetCommandLineA � EncodePointer �HeapAlloc GetLastError  �HeapFree  IsProcessorFeaturePresent �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �InterlockedIncrement  GetModuleHandleW  sSetLastError  �InterlockedDecrement  EGetProcAddress  �Sleep ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW WideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �HeapSize  %WriteFile GetModuleFileNameW  �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter  IsDebuggerPresent �RaiseException  9LeaveCriticalSection  � EnterCriticalSection  RtlUnwind rGetCPInfo hGetACP  7GetOEMCP  
IsValidCodePage �HeapReAlloc ?LoadLibraryW  -LCMapStringW  gMultiByteToWideChar iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  $WriteConsoleW � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll      �pQ    r          h l p ��    myplugin.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                         ��    .?AVNodeData@@  ��    .?AVBaseData@@  ��    .?AVObjectData@@    ��    .?AVContainerObject@@   ��    .?AVGeDialog@@  ��    .?AVGeModalDialog@@ ��    .?AVGeUserArea@@    ��    .?AVSubDialog@@ ��    .?AViCustomGui@@    ��    .?AVNeighbor@@  ��    .?AVC4DThread@@ ��    .?AVtype_info@@ u�  s�  cos             asin            sqrt            N�@���D        /a/a/a/a/a/a/a/a/a/a�������������
                                                                                           	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 ?         x�   |�   l�   p�   ��   ��!   ��   d�   \�   L�   ��   ��   0�   ,�    (�   D�   <�   ��   4�   ��   ��   ��   ��   ��"   ��#   ��$   ��%   ��&   ��      �      ���������              �       �D        � 0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     �%�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����C   ���������xl`XLHD@<840,($  �8������������	         xph`XPH8(������������|tl\H<0�$� � � � � � � p \                                                                                            �*            �*            �*            �*            �*                              h-        �(
��*`,    �&  8(     �            .   .   `-d@d@d@d@d@d@d@d@d@d-h@h@h@h@h@h@h@h-���   ���5      @   �  �   ����             �@    �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
    ����                                                                                                                                                                               �   0A0R0�0�0�0$181K1d1w1�1�1�1�112Q2b2�2�2�2�2�2�2A3Q3a3q3�3�3�3#434G4\4o4�4�4�45b5�5�6�6�6�6�6�6�6�6�6�6�6	7717E7X7t7�7�7�7�7�7	8888�8�89(9Q9�9�9 :B:l:�:;+;�;�;�;�;<B>I>f>�>D?�?�?    t   \0�0111G1d1x1�1�1K2`2�2k3�3�3j45 5�5
667@7V8$:�:�:�:-;];�;�;<<�<�<!=Q=}=�=�=�=>H>h>�>�>�>?T?�?�?�?   0  �   0H0m0�0�0�0!1T1�1�1�12I2�2�2383T3}3�3�3�3444b4�4�4�45-5a5�56-6a6�6�67-7]7�7�7�7H8h8�8�8�8949`9�9�9�9�9-:<<&<0<:<D<N<X<b<l<v<�<�<�<�<�<�<�=�?   @  \   	0/0]0�0�0�01�1�1�1&2L2�2�2�23B3i3�3�3�3�3(4X4�4�4�455O5s5�5�5�56�6�;l=p=t=x=|=   P  <   |2�2�2�2�2(353B3O3\3i3v3�3�3�3�3�<F=�=�>?-?T?�?�?�? `  h   90�2�2�2H344[4�4�4�45;5x5�5�5 6]6�6�6�6)7Y7�7�7�718m8�8	949a9�9�9�9�9!:T:�:�:�:�:/=�>�>)?Q?}?�? p  L   �4�4^5�5$6K6�6�6�67$7D7d7�7�78T8�8�8�819]9�9�9�9 :`:�:�:;�;<O?�? �  P   2%2+2q2�23L3b3�3�3�324r4�45Q5�5�56�6�67c7�78E8�8�89><>�>�>?y?�? �  8   #0s0/1G2�7`9�9�9�:3;�;�;=<�<�<S=�=>i>�>3?�?�?   �  p   R0�01r1�132�2�2C3�34�4"5h5�5�556w6�6�607s7�7#8c8�8�8�849�9�9:i:�:A;�;�;1<|<�<�<#=b=�=�=&>h>�>�>F?|?�? �  �   t0�0�2�3�3�3�3�3�3�3�3�3�355 5$5(5,50545856L6b6�6�6�67P7�7�7�78a8�8�8H9s9�9�9:Q:�:�:;3;l;�;�;=C=x=�=�=>H>x>�>�>0?i?{?�? �  T   00(0_0�0�0 1P1�1�1282h2�2�2S3�3�34@4o56E7�89�9�9:�:;\;y;=�=�=(>P>   �      B3�3�3#4$:(<<>�>�?�?�?   �  P   �0�2F3�3�3�3!4Q4�4�4�4�5�5�6�6�7�7�78M8H9h9�9�:%>U>m>�>�>�>?=?q?�?�?�? �  x   0C0�0�0�0m1�1�1�12Q2�2�2�213a3�3�3�3494i4�4�4�45=5t5�5�56(6H6h6�6�6�67M7}7�7�78=8m8H<W<�=�=�>�>?>?m?�?�?   �   010_0�0�0191T1x1�1�1�132h2�2�2�23(3H3h3�3�3�3 4P4y4�4�4�45=5]5�5i6�6�6�6	707\7�7�788�8�8 9P9�9�9�9	:(:H:m:�:�:�:-;];�;�;�;<M<}<�<�<===m=�=�=�=->a>�>�>�>)?t?�?�?  �   0>0n0�0�0111a1�1�1�12M2}2�2�23=3m3�3�34A4y4�4�45=5m5�5�5�5!6H6h6�6�6�67M7�7�7�7�8�89A9t9�9�9:/:c:�:�:�:#;T;�;�;�;�<�<=4=a=�=�=�=>M>}>�>�>?]?�?�?�?     \   !0Q0�0�0�0!1�1T2�2�2	363]3�3�3�3-4�4�4�45M5}5�56A6v6�6�67=7�7�7�7+8�9	:H:Z:�:�:> 0 L   22J2[2�4�4�4�4�6�6-7]7�7�7�7,8\8h8�8�89�9�9�9A:p:�:�=>Y>y?�?�?�? @ h   �0�01;1m1�1�1�12M2�2�23-3i3�3�3414t4�4�485]5�5�5�5$6M6�6�67d7�8�8989a9�9�9/:�:�:�:A;g>W?   P    w02�4�869   ` X   d6�7�7=8u8�8�8$9L99�9!:Q:=;o;�;�;�;-<d<�<�<�<=4=[=�=�=�=>P>�>�>�>)?`?�?�?�?   p �   %0M0}0�0�0�011d1�1�1�1�1 2M2i2�2�2�23N3y3�3�3�3	4)4I4d4�4�4�4�4	505Y5�5�5�56M6}6�6�67-7Y7�7�7�78@8�8�8 909`9�9�9�9:M:y:�:�:�:+;k;�;�;5<�<�<�<$=]=�=�=�=	>)>D>d>�>�>�>�>)?X? � �   090c0�0�0191Y1�1�12\2�2�2�2�2,3l3606l6�6�6�6 707`7�7�7�78D8p8�8�8�89@9p9�9�9�9:I:i:�:�:�:�: ;u;�;�;A<y<�<�<�<==y=�=�=!>D>s>�>�>$?T?�?�?�? � �   0Y0�0�0:1|1�1�1H2�2 3�3�34D4�45d5�5�5�56D6o6�6�67$7K7�7�7�78=8]8�8�8�89M9m9�9�9�9=:_:�:�:�:!;Q;�;�;�;<M<�<�<�<=3=c=�=   � 8   -2h2�2:Y;y;�;�;�;	<J<l<�<�<!=M=m=�=�=>->Y>o?�? � �   0-0Q0}0�0�0
1111J12I2�2�2�23A3q3�3�3-4�5�5�5$6D6q6�6�6�647]7�7�748�8�89d9�9�9�9�9�9�9:�:�:�:@;v;8<H<l<|<=�=|>�>�>�>�>�>?G?}?�?�?   � �   	0$0I0�0�0(1T1]1b1p1�1�1X2~2�2�2�2/3�3�3444"4[4b4�4�4�4�4�4�45.5D5H5L5P5T5X5m5�5�5�5#6s6�6717a7�7�7�7$8K8k8�8�8�89>9[9�9�9�9�9+:K:{:�:;+;[;{;�;<=<]<}<�<�<�<�<===]=}=�=�=�=�=>=>   � (   Z0i0�0�0s1�1�1�1�2�2�2�213F3D;   �    �;4<8<<<@<D<!>[>�?   � �   �12=2]2�2�2�2313d3�3�3414a4�4�4�4�6777777 7$7*7.73797=7C7G7M7Q7W7[7�7�7.8f8k8u8�8�8�8�89?9E9K9`9�9�9�9:F:�:�:�:1;6;?;N;q;v;{;�;<|<�<�<�<==(=B=�=�=�=	>>A>L>^>r>�>3?E?k?�?�?�?   �    00R0]0o0�0�0�0�0111191_1}1�1�1�1�1�1�1�1�1�1�1�1�1�1b2m2�2�2�2�2�2�2�23 3$3(3,3034383<3�3�3�3�3�3�3:4S4�4�4�45J5|5�5�5�5�5�5�5�5�56$6(6,6064686<6@6�6�6�6�6�677(7/74787<7]7�7�7�7�7�7�7�7�7�7�7&8,8084888�8�8Q9[9t9z9�9�9�9�:�:�:�:�=�=<>  $  �3]4�5�5 6;6@6K6R6^6d6p6v66�6�6�6�6�6�6�6�6�6�6�6�6	77D7�7�7�7�7�7�7�78�8�8�8�8�8G9W9]9i9o99�9�9�9�9�9�9�9�9�9�9�9�9�9�9:
::: :,:1:6:<:@:F:K:Q:V:e:{:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;C;L;X;�;�;�;�;�;�;<<<$<F<�<�<�<�<�<�<==#=-=C=N=h=s={=�=�=�=�=�=>>,>3>^>�>?	?3?x??�?�?�?     �   0(0F0j0�0�0�0�01181]1h1w1�1�1�122 2+2�3�34
444�4�4�4�45#52575X5]5�5�5�5�5�5�5�5"6�67777�7959B9N9V9^9j9�9�9�9�9�:�:�:
;";,;G;O;U;c;�;�;�;�;<S<�<�<�<�<�<3=@=F=e=j=�=�=�=�=�=>>>>�>�>?Y?�? 0 �   h0�0;1<2L2]2e2u2�233&3�3�3�3�3�3U4f4�4�4�4�4�4�4i5u5}5�5�56C6r6z6�6�6�7�7�7�9�9�9�9:C:|:�:�:�:�:�:�:�:;;H;c;j;s;|;�;�;�;�;�;�;�;<<<<<<#<'<+</<3<7<;<P<�<#=)=/=5=;=A=H=O=V=]=d=k=r=z=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>   @ �   1r2�2�2�2�2.374�4�4=5�5�7�7�7�7�7818t8�8%9�9�9�9�9�9:�:;';6;E;W;7<A<N<�<�<�<�<�<�<�< ==%=+=N=U=n=�=�=�=�=�=>\>|>�?�?   P �   �0o1�1�133D3~3�3�3�3�3�3�3�3�34"454Y4�4�4�4H5e5�56<6�6�6�6�6�677$7=7Y7b7h7q7v7�7�7�7�7�7F8�8�819�9":�:�:�:�:�;�;�<�<�=�? ` �   �1�1�1T2Z2f2�2�2�2 33333#3(383g3m3u3�3�3�3 44444&4�4�4�45�5�5�5�566�677$74797J7R7X7b7h7r7x7�7�7�7�7�7�7�7�78(8*:1:7:p:d;�;�<�<�=_>}>�>??-?   p @   {2k3�4�4%5F5&7G9K9O9S9W9[9_9c9<:�:�:%;?;H;p;�;R<"=�=�=X> � d   C2U2g2y2�2�2�2�2�2�233/3A3S3e3w3�3�4(56$6�6�7N8T8�8�8	9�9�9�9y:m;u;&<=�=�=F>L>Z>�>?G?�? � 4   �2�2�5�5�5�5�5�566
6666#6�677:7�7�7   � p   �1�3�3�3�34>4�405�5�5�67e7�8�9}:�:�:;$;�;�;<�<�< =2=8=R=a=n=z=�=�=�=�=�=�=�=�=>>B>u>�>�>�>�>??   � x   ,0J0W3j3�3�3�3464R44�4�4�4�455-5�5C6�6�6�6�6�677�788;8�8999$959�9:H:h:�:�:x;�;�;�; <2<Z<�<==&=D=   �   1111 1$1(14181�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2�2�2�5�5�5�5�5�5�5�5�5�566 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6X8\8`8�9�9�9�9�9�:�:�:`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�; � 4   <5D5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5�5�5�5 � �   �8�8�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   �    00000000 0$0(0,0004080<0@0D0H0L0P0T0X0�=�=>>>>4>8>P>`>d>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>??? ?0?4?<?T?d?h?x?|?�?�?�?�?�?�?�?�?�?�?�?  �   000040D0H0X0\0`0d0l0�0�0�0�0�0�0�0�0�0�0�0�01$1(181<1D1\1�1�1�1�1�12$2@2L2h2�2�2�2�2�23$3(3H3d3h3�3�3�3�34404P4p4     h   0000L0l0�0�0�0�0�01 1�1�1�1�1�1�1�1�1�1�1l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444$4,444<4D4L4�9�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<�<�<�<�<�<=(=,=0=4=8=D=H=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          