MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$       �]nQ�< �< �< {K��< �<�< v���< ���< v���< v���< v���< ���< ���< ���< Rich�<                         PE  L ���Q        � !  �  Z      q�                               p         @                   @2 O   �. <                            P �                                   @              �                           .text   %�     �                   `.rdata  �2      4   �             @  @.data   �   @                   @  �.reloc  "   P      "             @  B                                                                                                                                                                                                                                                                                                                                                                        �+  �   �����������������������L$t�   ùPA�  ������������  �����������VW�|$3���tfS�\$U�l$U�t$���NL  �|A�ϋ��   �@4�Ѕ�t��tj SU�t$$P�������|$$ t��|A�ϋ��   F�R(�ҋ���u�][_��^����������VW�|$3���tGS�\$U�l$���$    ��t$���K  ;�uF��u�|A�ϋ��   �@(�Ћ���u�][_��^�_��^���������j�h(�d�    P��$V�8A3�P�D$,d�    �|A�L$�@Q�@�С|Aj �@j��@�L$h� Q�Ѓ��D$P�L$�D$8    �fR  �|A�L$�@Q�@�D$8�С|A�L$ �@Q�@�С|Aj �@j��@�L$,h� Q�Ѓ�j �t$�D$$Ph� j j �D$L�  ��PhD� �3 �|A���I�D$8�IP�D$T�у� �L$�D$4�����S  �ƋL$,d�    Y^��0��̡|AQ�@�@��Y��t$��  Y������V����!  �D$t	V�  ����^� ��j�hi�d�    PQV�8A3�P�D$d�    jh�jEj��
  �����t$�D$    ��t ���R!  �4�ƋL$d�    Y^���3��L$d�    Y^���������SV�t$W�t$ ���t$ �t$ �t$ V�O  �؅�u_^[� ���> t	V��Z  ���O�LV  _�^��[� ��V�t$���N  ���> t	V�Z  ��^� ��������������̃�SV�t$$WV���>N  ����u	_^[��� �|AV�@@�@,�Ћ|A���Q���R4jh�  �������|A�D$���D$���D$�@�L$�@HQh�  ���Ѓ��; t	S�Z  ����_^[��� ������j�hq�d�    P��VW�8A3�P�D$ d�    �t$4�D$    �|A�L$�@Q�@(�Ћ��|A�|$8�IW�I�D$4   �ѡ|AW�@V�@�Ћ|A�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� �����������S�\$U�l$V�t$WUVS���M  �D$��u_^][� ��t4��t���F u4US���  �D$_^][� S���Y  �D$_^][� US���   �D$_^][� ����������j�h��d�    P��XSVW�8A3�P�D$hd�    ���L$|�?( �L$|HP�% � /������N  �$�  �t$xj jjj?���*�  P�t�������  �s�t$x3�Wjjj?����  P�Q�����  �R�|A�t$x���   �΋@4��j jjj?P�&������%�|A�t$x���   3��@4Wjjj?����P�������  �|A���@@V�@,�Ћ��D$$WP�������P�|AS�A�΋@8�D$x   �С|A�L$ �@Q�@�D$t�������U  �L$0�E  �D$LjP�D$x    �B  ��P�L$4�D$t�_%  �L$L�D$p �!  �|A�L$�@Q�@�Ѓ��D$Pj�D$x��
  ���L$4Pj j�Z!  �|A���I�D$�IP�D$t �у�����   �O����u	��V  ���R  ���uj�
  P�J�  ���Wj j��D$8P�7S  ��tj�;�  W�V  ���2�{V  j j��j@j@���*S  �jjh   V�S  W�cV  ���7�L$0�D$p�����   �L$hd�    Y_^[��d� � �Gt	P�)V  ���L$hd�    Y_^[��d� � . 
 � � 
 
 � � �����������̃�X�ISUVW�|$p��\$4�3��tL��tV�|Q  ��%Q  ���|AV�I�D$     �I�D$$    �ы|AV�I��I�D$�у��L��u�aU  j j��j@j@���R  ShD� ��3 ����t�V�Q  �C�k�D$�C�D$ �C�l$�D$����  �|A�t$l�@@�@,�Ћ|A���Q�����   j h�  ���҉D$$���  �|AW��L$8Q�D$<�D$D�D$L�@h�  ���   �L$XQ�����~ ���~P�~X�Y��Y��Y��,��ΉD$0�,D$,�,ÉD$(��R  �|A�؋ř����   �L$l�R4���D$$�D$�ҋ�����   j?���B  ��t�|A�ϋ��   �@(�Ћ���u��x   3�9l$~p�D$�L$��|^�|$ O|$�D$$�t$(�|A�t$0�@�t$8��  WUV�Ѓ���t�|Ah�   �@W��  USV�Ѓ�O�L$$u��D$�L$E;�|��L$l�^�  ������   �d$ j?����A  ��t�|A�ϋ��   �@(�Ћ���u��}   3�9l$~u�D$�L$��I ��|^�|$O|$�D$l�t$(�|A�t$0�@�t$8��  UWV�Ѓ���t�|Ah�   �@U��  WSV�Ѓ�O�L$lu��D$�L$E;�|��\$4�D$�C�D$ �C�D$�C�D$_�3�C�D$l^]�@   [��X� �G    _^][��X� j�h��d�    P�� VW�8A3�P�D$,d�    �|A�t$<�@@V�@,�Ѓ���j jj?����  P�����P�D$ P�F�����P�|Ah�  �A�ϋ@8�D$<    �С|A�L$�@Q�@�D$8�����С|A�����   �΋@4��j jj?P�z���P�D$0P�������P�|Ah�  �A�ϋ@8�D$<   �С|A�L$�@Q�@�D$8�����Ѓ��L$,d�    Y_^��,� �������������SVW�t$�|$W�t$���)E  �؅�u_^3�[� �D$P���4  ��t�N��t�M  ��Q  �F�|$ t�v���45  ��t�_^��[� ��������SVW�|$W�t$����D  ��3���t89F����P�w2  ��u_^3�[� �F��tjj h�� P����2  ��t܋�_^[� ������̋|A�D$��t<�|$ �t$�I�t$�   t;�B�P���   �Ѓ�Ã�B�P���  �Ѓ�ù   ;�VB�W�xW�� ������u_^À|$ tWj V輵 �������_�F�LA   ^�����������̋L$��t,�=LA t�y���A�u
�D$�%� �|A�L$�@� �������������̋L$��t�|A�L$�@��@  �����̡|Ahﾭދ@��@  ��Y����������V�t$���t�|AQ�@� �Ѓ��    ^�������������̡|A�@���  ���D$��t�x��u�   �3����������̡|A�@��  ��|A�@��   ���D$�   ;�VB�W�xW�� ������u_^Ã|$ tWj V�b� �������_�F�LA   ^���    �A    �A    �A    �����V��~ u=���t�|AQ�@<�@�Ѓ��    W�~��t���  W�U������F    _^���������j�h�d�    P��V�8A3�P�D$$d�    ��D$P��7  ��P���D$0    �-   �L$���D$,�����  �ƋL$$d�    Y^��(��������j�h<�d�    PQV�8A3�P�D$d�    ��~ uTjh�j;j��������D$�D$    ��t�t$���  �3��D$�����F��u�L$d�    Y^��� �~ t3�9�"�|A�t$�@<� �Ћȃ�3���F   �����L$d�    Y^��� ��������������V���F   �|A�@<�@��3Ʌ����^��������������̋	�|A��u�@� � �@<�t$�@Q�Ѓ�� ���������̃y t�   ËQ��u3�á|AR�@<�1�@�Ѓ��������V��~ u=���t�|AQ�@<�@�Ѓ��    W�~��t����  W�5������F    _^��������̋PA�|A��u�@� Ë@<�t$�@Q�Ѓ������������j�h��d�    P��(SV�8A3�P�D$4d�    �D$    �PA��u�|A�A�0��|A�t$H�@<Q�@�Ћ|A�����I�D$�IP�ѡ|A�L$�@Q�@V�С|A�L$0�@Q�@�D$L   �С|Aj �@j��@�L$<h@Q�Ѓ� �|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@��tA�t$D�@V�Ћ|A�D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С|Aj��@j��t$T�@L�t$�L$$�С|A�t$D�@V�@�С|A�L$�@V�@Q�Ћ|A�D$ �IP�I�D$    �D$L �у��ƋL$4d�    Y^[��4��j�h��d�    P��(SV�8A3�P�D$4d�    �D$    �PA��u�|A�A�0��|A�t$H�@<Q�@�Ћ|A�����I�D$�IP�ѡ|A�L$�@Q�@V�С|A�L$0�@Q�@�D$L   �С|Aj �@j��@�L$<hDQ�Ѓ� �|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@��tA�t$D�@V�Ћ|A�D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С|Aj��@j��t$T�@L�t$�L$$�С|A�L$$�@Q�@�С|Aj �@j��@�L$0hHQ�Ѓ��|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@��t�t$D�@V�������@Hj�t$�L$�С|Aj��@j��t$X�@L�t$�L$$�С|A�t$D�@V�@�С|A�L$�@V�@Q�Ћ|A�D$ �IP�I�D$    �D$L �у��ƋL$4d�    Y^[��4����������j�h �d�    P��(SV�8A3�P�D$4d�    �D$    �PA��u�|A�A�0��|A�t$H�@<Q�@�Ћ|A�����I�D$�IP�ѡ|A�L$�@Q�@V�С|A�L$0�@Q�@�D$L   �С|Aj �@j��@�L$<hLQ�Ѓ� �|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@��tA�t$D�@V�Ћ|A�D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С|Aj��@j��t$T�@L�t$�L$$�С|A�L$$�@Q�@�С|Aj �@j��@�L$0hPQ�Ѓ��|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@��t�t$D�@V�������@Hj�t$�L$�С|Aj��@j��t$X�@L�t$�L$$�С|A�L$$�@Q�@�С|Aj �@j��@�L$0hTQ�Ѓ��|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@���D����@Hj�t$�L$�С|Aj��@j��t$\�@L�t$�L$$�С|A�t$D�@V�@�С|A�L$�@V�@Q�Ћ|A�D$ �IP�I�D$    �\$L�у��ƋL$4d�    Y^[��4��������������j�h|�d�    P��(SV�8A3�P�D$4d�    �D$    �PA��u�|A�A�0��|A�t$H�@<Q�@�Ћ|A�����I�D$�IP�ѡ|A�L$�@Q�@V�С|A�L$0�@Q�@�D$L   �С|Aj �@j��@�L$<hXQ�Ѓ� �|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@��tA�t$D�@V�Ћ|A�D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С|Aj��@j��t$T�@L�t$�L$$�С|A�L$$�@Q�@�С|Aj �@j��@�L$0h\Q�Ѓ��|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@��t�t$D�@V�������@Hj�t$�L$�С|Aj��@j��t$X�@L�t$�L$$�С|A�L$$�@Q�@�С|Aj �@j��@�L$0h`Q�Ѓ��|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@���D����@Hj�t$�L$�С|Aj��@j��t$\�@L�t$�L$$�С|A�L$$�@Q�@�С|Aj �@j��@�L$0hdQ�Ѓ��|Aj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ��|A�L$$�@Q�@���D$@�С|A���@��������@Hj�t$�L$�С|Aj��@j��t$`�@L�t$�L$$�С|A�t$D�@V�@�С|A�L$�@V�@Q�Ћ|A�D$ �IP�I�D$    �\$L�у��ƋL$4d�    Y^[��4ËD$�PA��EȉL$� �������̡|A�@<�@����̋D$����u���VP�L$� �D$P�D$P�L$�D$    �D$    �� ����   �t$��$    �D$��tB��t=��uZ�|A�t$���   �@H�Ћ|A�ЋA���@xV���Ѕ�u,�   ^��á|A�t$���   �@T��VP�J�������uԍD$P�D$P�L$�@ ���x���3�^����j�h��d�    P��HSUVW�8A3�P�D$\d�    3ۉ\$�|A�L$,�@Q�@�С|AS�@j��@�L$8hhQ�С|A�L$@�@<Q�@�\$|�Ћ|A���I�D$D�IPǄ$�   �����у���u3��L$\d�    Y_^][��T�V�L$(3��( �D$P�D$$P�L$,�e ���  �l$l���$    �|$ ��   �|A�t$���   �@T�Ћ�����tc�|A�D$<�IP�I�у��D$<Pj�D$T��P���D$p   �\$$�p  �Ћ|A���AU�@x���D$h   �\$���D$��t�D$ �D$d   ��t�|A�L$L�@����@Q�\$�Ѓ��D$d������t�|A�L$<�@Q�@����Ѓ��|$ u�D$P�D$$P�L$,�X ��� �����|$�ǋL$\d�    Y_^][��T�����j�h&�d�    P��DSUVW�8A3�P�D$Xd�    �t$l3ۉ\$��u|�|A�L$(�@Q�@�С|AV�@j��@�L$4htQ�С|A�L$<�@<Q�@�t$x�Ћ|A���I�D$@�IP�D$|�����у���u3��L$Xd�    Y_^][��P�V�L$$3��# �D$P�D$ P�L$(�` ����   �|$h�d$ �D$����   �|A�t$���   �@T�Ћ�����tc�|A�D$8�IP�I�у��D$8Pj�D$P��P���D$l   �\$$�n  �Ћ|A���AW�@x���D$d   �\$���D$l��t�D$l �D$`   ��t�|A�L$H�@����@Q�\$�Ѓ��D$`������t�|A�L$8�@Q�@����Ѓ��|$l tR�l$�ŋL$Xd�    Y_^][��PÃ�u3�L$��t+�|AQ���   �@H�Ћ|A�ЋA���@xW���Ѕ�t��D$P�D$ P�L$(� �����������������̡|A�@<�@����̃=XA uK�PA��t�|AQ�@<�@�Ѓ��PA    V�5\A��t���  V��������\A    ^������������j�hq�d�    P��VW�8A3�P�D$ d�    �t$8�D$    �|A�t$8�@�T$���   R�Ћ��|A�|$0�IW�I�D$,   �ѡ|AW�@V�@�Ћ|A�D$�IP�I�D$   �D$8 �у��ǋL$ d�    Y_^�� � ������������������������̅�t�j������̡|A�@��  ��|A�@��(  ��j�h��d�    P�� �8A3�P�D$$d�    �D$    �|A�T$�@R��   �ЋL$4P�D$0   �  �L$�D$   �D$, �  �D$4�L$$d�    Y��,� �̡|A�@��$  ��|A�@��  ��|A�@���  ��|A�@��  ��|A�@���  ��|A�@��x  ��|A�@��|  ��|A�@��d  ��|A�@��p  ��|A�@��t  ���D$V����t	V�z�������^� ̡|A�@$�@X����̡|A�@$�@\������t$�|A�t$�@$�t$�@`Q�Ѓ�� j�h��d�    PQV�8A3�P�D$d�    ��t$�|AV�@�@�С|AV�@$�D$    �@D�Ѓ��ƋL$d�    Y^�����������������j�h��d�    PQV�8A3�P�D$d�    ��t$�|AV�@�@�С|AV�@$�D$    �@D�С|A�t$$�@$V�@d�Ѓ��ƋL$d�    Y^��� ����������j�h�d�    PQV�8A3�P�D$d�    ��t$�|AV�@�@�С|AV�@$�D$    �@D�С|A�t$$�@$V�@�Ѓ��ƋL$d�    Y^��� ����������j�hA�d�    PQV�8A3�P�D$d�    ��t$�|AV�@�@�С|AV�@$�D$    �@D�С|AV�@$�t$(�@L�Ѓ��ƋL$d�    Y^��� ����������j�hd�d�    PQV�8A3�P�D$d�    ��t$�|AV�@$�D$    �@H�С|AV�@�D$�����@�Ѓ��L$d�    Y^����������̡|A�t$�@$Q�@L�Ѓ�� �������̡|A�@$�@����̡|AQ�@$�@�Ѓ����������������j�h��d�    P��VW�8A3�P�D$ d�    �D$    �|AQ�@$�L$�@Q�Ћ��|A�|$8�IW�I�D$4   �ѡ|AW�@V�@�Ћ|A�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� � ����������̡|A�t$�@$Q�@�Ѓ�� ��������j�h��d�    P�� VW�8A3�P�D$,d�    �D$    �|AQ�@$�L$�@ Q�Ћ��|A�|$D�IW�I�D$@   �ѡ|AW�@$�D$D�@D�С|AW�@$V�@L���D$$   �|A�L$(�@$Q�@H�D$P   �Ћ|A�D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,� ��������������j�h8�d�    P�� VW�8A3�P�D$,d�    �D$    �|AQ�@$�L$�@$Q�Ћ��|A�|$D�IW�I�D$@   �ѡ|AW�@$�D$D�@D�С|AW�@$V�@L���D$$   �|A�L$(�@$Q�@H�D$P   �Ћ|A�D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,� ��������������j�h|�d�    P�� �8A3�P�D$$d�    �D$P�D$    ������t$4���D$0   �(����D$   �|A�L$�@$Q�@H�D$0   �Ћ|A�D$�IP�I�D$4 �ыD$<���L$$d�    Y��,� ����̡|AQ�@$�@(��Yá|AQ�@$�@h��Yá|A�t$�@$Q�@,�Ѓ�� �������̡|A�t$�@$Q�@0�Ѓ�� �������̡|A�t$�@$Q�@4�Ѓ�� �������̡|A�t$�@$Q�@8�Ѓ�� �������̡|A�t$�@$�t$�@PQ�Ѓ�� ���̡|A�t$�@$Q�@T�Ѓ�� �������̡|A�@$�@l����̡|A�@$�@p����̡|AV�@$��@LV�t$�Ѓ���^� ��j�h��d�    PQV�8A3�P�D$d�    �D$    �|A�t$�@V�@�D$    �С|AV�@$�D$   �@D�С|AV�@$�t$,�@L�Ћ|A�t$4�I$V�I@�D$,    �D$    �у��ƋL$d�    Y^�������������̡|AV�@$�t$�@@��V�Ѓ���^� �̡|A�t$�@$Q�@<�Ѓ�� �������̡|A�t$�@$Q�@<�Ѓ����@� ���j�h��d�    P��VW�8A3�P�D$ d�    �D$    �|AQ�@$�L$�@tQ�Ћ��|A�|$8�IW�I�D$4   �ѡ|AW�@V�@�Ћ|A�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� � ����������̡|A�@(�@����̡|A�@(�@����̡|A�@(�@����̡|A�@(�@����̡|A�@(�@ ����̡|Aj�t$�@(�t$�@��� �������t$�|A�t$�@(�t$�@$��� ���̡|A�@(�@(����̡|A�@(�@,����̡|A�@(�@0����̡|A�@(�@4����̡|A�@(�@X����̡|A�@(�@\����̡|A�@(�@`����̡|A�@(�@d����̡|A�@(�@h����̡|A�@(�@l����̡|A�@(�@p����̡|A�@(�@t����̡|A�@(�@x����̡|A�@(���   ��j�h�d�    P��V�8A3�P�D$d�    ��|A�L$�@Q�@�Ѓ��D$P���D$$    �   ��u3���|A�L$�@$Q�t$,�@�Ѓ��   �|A�D$�IP�I�D$$�����у��ƋL$d�    Y^��� ��������Q�|A�T$�@(R�@X�Ѕ�uY� �D$3�8L$����   Y� �������������j�h:�d�    P��V�8A3�P�D$ d�    ��|A�D$    �D$    �@(�L$�@hQ���Ѕ���   �L$�|A��uM�@�L$�@Q�С|A�t$4�@�L$�@Q�D$4    �С|A�L$�@Q�@�D$8�����Ѓ��   �@h����   hj  Q�Ћȡ|A���L$�@(��u�@4j�����3��L$ d�    Y^��$� �@j �t$Q���Ѕ�u"�D$P������3��L$ d�    Y^��$� �|Aj �H�D$HP�t$�A�t$<�ЍD$P�@������   �L$ d�    Y^��$� ����̡|AV�@(W�|$�@pW���Ѕ�t8�|A�΋P(�GP�Bp�Ѕ�t!�|A�΋P(�GP�Bp�Ѕ�t
_�   ^� _3�^� ������̡|AV�@(W�|$�@tW���Ѕ�t8�|A�΋P(�GP�Bt�Ѕ�t!�|A�΋P(�GP�Bt�Ѕ�t
_�   ^� _3�^� ������̡|AS�@(V�@pW�|$W���Ѕ���   �|A�΋P(�GP�Bp�Ѕ���   �|A�΋P(�GP�Bp�Ѕ�tn�|A�_�@(S�@p���Ѕ�tW�|A�΋P(�CP�Bp�Ѕ�t@�|A�΋P(�CP�Bp�Ѕ�t)�GP��������t�G$P��������t_^�   [� _^3�[� ��������̡|AS�@(V�@tW�|$W���Ѕ���   �|A�΋P(�GP�Bt�Ѕ���   �|A�΋P(�GP�Bt�Ѕ�tn�|A�_�@(S�@t���Ѕ�tW�|A�΋P(�CP�Bt�Ѕ�t@�|A�΋P(�CP�Bt�Ѕ�t)�G0P���/�����t�GHP��� �����t_^�   [� _^3�[� ��������̡|A�@(�@8����̡|A�@(�@<����̡|A�@(�@@����̡|A�@(�@D����̡|A�@(�@H����̡|A�@(�@L����̡|A�D$�@(Q�@P�$��� ���̡|A�D$�@(���@T�$��� �̡|A�t$�@(�t$�@|��� �������̡|A�t$�@(�t$���   ��� �����j�h]�d�    P��V�8A3�P�D$d�    ��L$(�D$P����P���D$$    �\   �|A���I�D$�IP�D$$�����у��ƋL$d�    Y^��� ������̡|A�|$ �P(�����D$�B8������Q�|AV�@W�@d���L$j �Ћ|Ah��I�p���   h�  V�ыȡ|A���L$��u�@(j��@4����_3�^Y� �@j �@hVQ�L$�С|AV�@(�ϋ@H�Ѕ�t2�|AV�@(�t$�@ ���Ѕ�t�D$P�   ��������_^Y� �D$P3���������_^Y� �����̡|AV�@(W�|$�@P�Q���$�Ѕ�tF�|A�G�@(Q�@P���$�Ѕ�t(�|A�G�@(Q�@P���$�Ѕ�t
_�   ^� _3�^� �|AV�@(W�|$�@T������$�Ѕ�tJ�|A�G�@(���@T���$�Ѕ�t*�|A�G�@(���@T���$�Ѕ�t
_�   ^� _3�^� ���������̡|AV�@(W�|$�@P�Q���$�Ѕ��  �|A�G�@(Q�@P���$�Ѕ���   �|A�G�@(Q�@P���$�Ѕ���   �|A�G�@(Q�@P���$�Ѕ���   �|A�G�@(Q�@P���$�Ѕ���   �|A�G�@(Q�@P���$�Ѕ�ts�|A�G�@(Q�@P���$�Ѕ�tU�|A�G�@(Q�@P���$�Ѕ�t7�|A�G �@(Q�@P���$�Ѕ�t�G$P���������t
_�   ^� _3�^� ��������̡|AV�@(W�|$�@T������$�Ѕ���   �|A�G�@(���@T���$�Ѕ���   �|A�G�@(���@T���$�Ѕ���   �|A�G�@(���@T���$�Ѕ�th�|A�G �@(���@T���$�Ѕ�tH�|A�G(�@(���@T���$�Ѕ�t(�G0P���T�����t�GHP���E�����t
_�   ^� _3�^� �|A�@(� �����̡|AV�@(�t$�@�6�Ѓ��    ^�̡|A�@(���   ��|A�@(�@����̡|A�@(�@����̡|AV�@(�t$�@�6�Ѓ��    ^�̡|A�t$�@,�t$�@Q�Ѓ�� ���̡|A�@,�@����̡|A�@,�@����̡|A�@,�@����̡|A�@,�@ ����̡|A�@,�@(����̡|A�@,�@$����̡|A�@,�@�����j�h��d�    P�� VW�8A3�P�D$,d�    �D$    �|A�T$�@,R�@�Ћ��|A�|$<�IW�I�D$8   �ѡ|AW�@$�D$<�@D�С|AW�@$V�@L���D$   �|A�L$ �@$Q�@H�D$H   �Ћ|A�D$$�IP�I�D$L �у��ǋL$,d�    Y_^��,� ��������������̡|Aj �@,j � �Ѓ�������������̡|AV�@,�t$�@�6�Ѓ��    ^�̡|A�@,�@4����̡|A�@,�@8�����j�h��d�    P�� VW�8A3�P�D$,d�    �D$    �|A�T$�@,R�@<�Ћ��|A�|$<�IW�I�D$8   �ѡ|AW�@$�D$<�@D�С|AW�@$V�@L���D$   �|A�L$ �@$Q�@H�D$H   �Ћ|A�D$$�IP�I�D$L �у��ǋL$,d�    Y_^��,� ���������������j�h1�d�    P��VW�8A3�P�D$ d�    �t$4�D$    �|A�T$�@,R�@@�Ћ��|A�|$0�IW�I�D$,   �ѡ|AW�@V�@�Ћ|A�D$�IP�I�D$   �D$8 �у��ǋL$ d�    Y_^�� � �������̡|A�@,�@,����̡|AV�@,�t$�@0�6�Ѓ��    ^�̡|A�@���  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@�@����̡|A�@�@����̡|A�@�@����̡|A�@�@����̡|A�@�@����̡|A�@�@����̡|A�t$�@�t$�@\��� �������̡|A�t$�@�t$��  ��� ����̡|A�D$�@���@ �$��� �̡|A�D$�@Q�@$�$��� ���̡|A�D$�@���@(�$��� �̡|A�@�@,����̡|A�@�@0����̡|A�@�@4����̡|A�@�@8����̡|A�@�@<����̡|A�@�@@����̡|A�@�@D����̡|A�@�@H����̡|A�@�@L����̡|A�@�@P����̡|A�@���   ��|A�t$�@Q��  �Ѓ�� ����̡|A�@�@T����̡|A�@�@X����̋T$��u3�� �|AR�@ Q�@(�Ѓ��   � ��������̡|A�@���   ��|A�@�@`����̡|A�@�@d����̡|A�@�@h����̡|A�@�@l����̡|A�@�@p����̡|A�@�@t����̡|A�@���   ��|A�@��  ��|A�@�@x����̡|A�@�@|����̡|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�t$�@Q��  �Ѓ�� ����̡|A�@���   ��|A�@���   ���T$��t�|AR�@ Q�@$�Ѓ���t�   � 3�� ����̡|AQ�@ �t$�@L�t$�Ѓ�� ���̡|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|AV�@�t$���   V�Ѓ��    ^���������������̡|A�@� �����̡|A�@�@����̡|A�@���   ��|A�@��   ��|A�@�@����̡|A�@�@����̡|A�@�@����̡|A�@�@����̡|A�@�@����̡|A�@���  ��|A�@�@�����j�h\�d�    P��V�8A3�P�D$$d�    �t$4�D$P�������|A�L$�@$Q�@�D$0    �Ѓ���t_�|A�L$�@j�@Q�Ѓ���u�D$P��������t3�|Aj�@V�@�Ѓ���u�|AV�@�@�Ѓ���t�   �3��|A�L$�@$Q�@H�D$0   �Ћ|A�D$�IP�I�D$4�����у��ƋL$$d�    Y^��(���������������̡|A�@�@ ����̡|A�@�@(����̡|A�@��  ��|A�@��   ��|A�@��  ��|A�@��  ��j�h��d�    P�� VW�8A3�P�D$,d�    �D$    �|A�L$�@Q�@$�Ћ��|A�|$@�IW�I�D$<   �ѡ|AW�@$�D$@�@D�С|AW�@$V�@L���D$    �|A�L$$�@$Q�@H�D$L   �Ћ|A�D$(�IP�I�D$P �у��ǋL$,d�    Y_^��,��j�h��d�    P�� VW�8A3�P�D$,d�    �D$    �|A�L$�@Q���  �Ћ��|A�|$@�IW�I�D$<   �ѡ|AW�@$�D$@�@D�С|AW�@$V�@L���D$    �|A�L$$�@$Q�@H�D$L   �Ћ|A�D$(�IP�I�D$P �у��ǋL$,d�    Y_^��,���������������Qj�t$�D$    �  �D$�������j�hz�d�    P��<SVW�8A3�P�D$Ld�    �D$    ��A��t�D$0P�^������D$T   �   �@�|A�L$�@Q�@�С|A�L$�@$Q�@D�D$\   �Ѓ��|$�D$T   �   �|A�t$\�@V�@�\$�С|AV�@$�D$\   �@D�С|AV�@$W�@L�Ѓ�����t;����\$�|A�L$�@$Q�@H�D$X   �С|A�L$�@Q�@�D$\�Ѓ��D$T    ��t<����\$�|A�L$0�@$Q�@H�D$X   �Ћ|A�D$4�IP�I�D$\ �у��ƋL$Ld�    Y_^[��H���������������j�h��d�    P�� VW�8A3�P�D$,d�    �t$@�D$    �|A�L$�@Q���  �Ћ��|A�|$D�IW�I�D$@   �ѡ|AW�@$�D$D�@D�С|AW�@$V�@L���D$$   �|A�L$(�@$Q�@H�D$P   �Ћ|A�D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,����������̡|A�@��D  ��|A�@��H  ��|A�@��L  ��j�h�d�    P��VW�8A3�P�D$ d�    �t$8�D$    �|A�t$8�@�L$���  Q�Ћ��|A�|$<�IW�I�D$8   �ѡ|AW�@V�@�Ћ|A�D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� ���̡|A�@���  ��|A�@���  ���A    �    �A    �A   ������t$�|A�t$�@@�t$�@Q�Ѓ�� �|A�t$�@@Q�@�Ѓ�� �������̡|A�t$�@@�t$�@Q�Ѓ�� ���̡|A�t$�@@Q�@ �Ѓ�� �������̡|A���   �@��|A���   �@��|A���   �@ ��|A���   �@$��|A���   ���   ��������������̡|A���   ��D  ��������������̡|A�t$�@@Q�@L�Ѓ�� �������̡|AQ�@@�@H�Ѓ���������������̡|A���   ���   ��������������̡|A���   ���   ��������������̡|AQ�@H���   �Ѓ�������������V��L$��t2�T$�|A���   ��t
�@@R��^� �T$�@D��tR��^� V��^� ��������������̡|A�@@�@0�����V�t$���t�|AQ�@@�@�Ѓ��    ^������������̡|AV�@@��@V�ЋЋD$����t��#��С|AR�@@V�@�Ѓ�^� �����t$�D$�|A�����   �$�t$���   �t$�t$�t$��� �������̡|A���   ���   ��������������̡|AQ�@H���   �Ѓ������������̡|A�t$�@HQ��d  �Ѓ�� ����̡|A�@@�@T����̡|A�@@�@X����̡|A�@@�@\����̡|A�@@�@`����̡|A�@@�@d����̡|A�@@�@h����̡|A�@@�@l����̡|A�@@���   ��|A�@@�@t����̡|A�@@�@x����̡|A�@@�@|����̡|A�@@���   ��|A�@@���   ��|A�@@���   ��|A���   �@t��|A�@@���   ��|A�@@���   ��|A�@@���   ��|A�@@���   ��|A�@@���   ��|A�@@���   ��|A�@@���   ��V�t$���t�|AQ�@@�@�Ѓ��    ^������������̡|A�@@�@0����̡|Aj�@@�L$�@4Qj �Ѓ�������̡|Aj�@@�L$�@4Qh   @�Ѓ����̡|A�t$�@@�t$�@4j �Ѓ������̡|A�@|� ������V�t$���t�|AQ�@|�@�Ѓ��    ^������������̡|A�@|�@ �����V�t$���t�|AQ�@|�@(�Ѓ��    ^������������̡|A�@ �@H����́|$qF uKW�|$��tA�|A�t$���   �ϋ@D�С|A�t$�@@�@,�Ћ|A���ЋAW�t$�@p����_����������̡|A�@��T  ��|AS�@@V�@,W�t$�Ћ|A�t$�I@�؋I,�ы|A���yh��hE  �ˋ��	�  Ph��hE  �����  P��T  �Ѓ�_^[�������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������3�� �����������3�� ����������̋L$�D$�A4�D$�A �D$��D$�A0�D$�AP4 �A8�e �A<�e �A@f �AD�e �AH�e �AL�e �AP�e �Al�e �AX�e �A\�e �A`f �Ad�e �AT�e �Ah�e �Ap	f �Atf �A(�A,    �����������́�   h�   �D$j P�!p j ��$�   �D$��$�   ��$�   ��$�   P������$�   h�   �D$T�D$(P��$�   ��$�   j�7�  ���   �j�hV�d�    P��   SV�8A3�P��$�   d�    ����	  ����H  ��$�   �L$ �����|A�L$�@Q�@Ǆ$�       �С|Aj �@j��@�L$h�Q�Ѓ��D$P�L$<Ƅ$�   �S�����$�   PƄ$�   �.����L$<QP�D$|PƄ$�   �6����L$,QP�D$lPƄ$�   �������j j�PƄ$�   ��  ���L$T��Ƅ$�   ������L$pƄ$�   �������$�   Ƅ$�   �����L$8Ƅ$�   �����|A�L$�@Q�@Ƅ$�    �Ѓ��L$Ǆ$�   �����y�����t	V�  ���Ƌ�$�   d�    Y^[�Ĩ   � V�t$����  �����^� ���������Q�j  YË�`��`��`��`��`��`��` ��`$��`(��`,��`0��`4��`8��`<��`@��`�������̡|A�@��   ��|AV�@�t$��$  �6�Ѓ��    ^��������������̡|AV�@��(  V�t$�Ѓ���^� ��������������̡|AQ�@�t$��,  �Ѓ�� ����̡|AQ�@�t$��,  �Ѓ����@� �D$��t�P�3ҡ|AR�@Q��8  �Ѓ�� ��������̡|A�t$�@Q��<  �Ѓ�� ������t$�|A�t$�@�t$��@  Q�Ѓ�� ������������̡|A�t$�@�t$��D  Q�Ѓ�� ̡|A�t$�@Q��H  �Ѓ�� �����j�h��d�    P��VW�8A3�P�D$ d�    �t$4�D$    �|AQ�@�L$��L  Q�Ћ��|A�|$<�IW�I�D$8   �ѡ|AW�@V�@�Ћ|A�D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� � ���̡|AQ�@��T  �Ѓ������������̡|AQ�@��P  �Ѓ������������̡|A�t$�@Q��X  �Ѓ�� ����̡|A�t$�@Q��l  �Ѓ�� ����̡|A�@��0  ��|A�@��4  ��|A�@��p  ��|A�@��t  ��|A�@��\  ��|AV�@�t$��`  �6�Ѓ��    ^����������������t$�|A�t$�@�t$��d  �t$�t$Q�Ѓ�� ������t$�|A�t$�@�t$��h  �t$�t$Q�Ѓ�� ����̡|AQ�@�@�Ѓ�����������������t$�|A�t$�@�t$�@X�t$Q�Ѓ�� �����������̡|A�t$�@Q�@\�Ѓ�� �������̡|AQ�@�@ ��Y�j�h��d�    P��V�8A3�P�D$d�    �|Ah�  �@Q���   �L$Q��P�|A�D$0    ���   �@8�Ћ|A�����   �D$�	P�D$4�����у��ƋL$d�    Y^����̡|A�@��   ���t$�|A�t$�@�t$�@Q�Ѓ�� �t$�|A�t$�@�t$���   �t$Q�Ѓ�� ��������̡|A�@�@$������t$�|A�t$�@�t$�@(�t$Q�Ѓ�� �������������t$�|A�t$�@�t$�@,�t$Q�Ѓ�� �������������t$$�|A�t$$�@�t$$�@`�t$$�t$$�t$$�t$$�t$$�t$$Q�Ѓ�(�$ �������̡|AV�@W�@��W�Ћ|AW�J���I���t$�|A�t$�Q�t$�N�QHP�B4j j W�Ѓ�(_^� �t$�|A�t$�@�t$�@4�t$�t$�t$�t$Q�Ѓ� � �|A�t$�@�t$�@@Q�Ѓ�� ���̡|A�t$�@Q�@D�Ѓ�� �������̡|AQ�@�@L�Ѓ���������������̡|AQ�@�@L�Ѓ���������������̡|AQ�@�@P�Ѓ���������������̡|A�t$�@Q�@T�Ѓ�� �������̡|A�t$�@Q�@T�Ѓ�� �������̡|AQ�@�@h�Ѓ���������������̡|A�t$�@�t$���   Q�Ѓ�� �j�h �d�    P��V�8A3�P�D$d�    �t$4�D$    �|A�t$4�@Q���   �L$Q�ЋЋt$<j �    �F    �|AR���   V�@�D$@   �Ћ|A�D$(���   P�	�D$(   �D$D �у� �ƋL$d�    Y^�� � �����������̡|A�@� �����̡|AV�@�t$�@�6�Ѓ��    ^���t$�|A�t$�@�t$���   �t$�t$Q�Ѓ�� ����̡|AV�@�t$�@�6�Ѓ��    ^��QS�\$V�C    �|A��@V�@h�Ѓ����|Au �@h���0  h�  �Ѓ�^3�[Y� �L$Q�L$Q�t$�D$    �@V���   �Ѓ���t�3�9t$~+W�d$ �D$�<� �<�tj����  ��t��F;t$|�_�D$P�`������   ^[Y� ��QS�\$V�C    �|A��@V�@h�Ѓ����|Au �@h���0  h�  �Ѓ�^3�[Y� �L$Q�L$Q�t$�D$    �@V���   �Ѓ���tσ|$ t�3�9t$~?W�D$����t+�|AQ�@�@h�Ѓ���t�D$j�<����  ��t�8F;t$|�_�D$P腮�����   ^[Y� ������̡|A�@��x  ��|A�@��|  ��|AQ�@���   �Ѓ������������̡|A�t$�@Q���   �Ѓ�� ����̡|A�@���   ��|AV�@�t$���   �6�Ѓ��    ^���������������VW���O����W�f�G f�G(f�G0f�G8f�G@f�GHf�GPf�GX�    �G`    �Gd    �Gh    �Gp�Gx�����G|   ��_^�������j�h&�d�    PQV�8A3�P�D$d�    ��t$�D$    �k   �N�D$�����[����L$d�    Y^�������������W��    �A`    �Ad    �Ah    �Ap�Ax�����A|   ���������������SW�����t7���_����xP t$V���Q���j j �pPj�GP���=����H ���^�    �O`��t�|AQ�@�@�Ѓ��G`    _[��������������j�h]�d�    PQ�8A3�P�D$d�    jh(h�   h�   ��������D$�D$    ��t���/����L$d�    Y���3��L$d�    Y����������������j�h��d�    PVW�8A3�P�D$d�    �|$�7��t,�t$���D$    ������N�D$���������V��������    �L$d�    Y_^��á|AS�@U�l$��   VW��W�_dS�wx�w`UV�Ѓ��G|����   �? ��   �; ��   �wpV�_hSU��  ����u&�W���|Ahx�@h  ��0  �Ѓ��wU�������j j jV��  �G|��t��������G|_^][� �G|�Gx����_^][� �G|�����    �|A�6�@�@�Ѓ��    �G|_^][� �����������V������W��    �F`    �Fd    �Fh    �Fp�Fx�����F|   ^������W���d �G`t~S�\$;_xtsU�/�͉D$謿���xP u����%V��虿��S�t$�pPj�GP��脿���H ���^�G|]��u�D$�_x��t�    �G`[_� �L$�Gx������t�3�[_� �̋D$��t	�Ap� �yd t�Ah� 3��y|��� ��������t$�|A�t$�@�t$�@�t$�t$�t$�t$Q�Ѓ� � �|A�t$�@Q�@�Ѓ�� �������̡|AQ�@�@��Yá|A�t$�@�t$�@Q�Ѓ�� ���̡|A�@� �����̡|AV�@�t$�@�6�Ѓ��    ^��VW���W����t$���t$�x@�t$�A����H ���_^� �����VW���'����t$���t$�xD�t$�����H ���_^� �����W��������xH u3�_�V�������ύpH�ܽ���H �^_�����W���Ƚ���xL u3�_� V��贽���t$���t$�pL�t$螽���H ���^_� ��W��舽���xP u���_� V���s����t$���t$�pP�t$�t$�Y����H ���^_� �������������W���8����xT u���_� V���#����t$���t$�pT�����H ���^_� �����W��������xX u���_� V�������t$�ύpX�ռ���H ���^_� ���������j�h��d�    P��$SVW�8A3�P�D$4d�    �ً|$D��tA�L$ ��  ���D$<    �x����pL�D$ P���i����H ��ЍL$ ��D$<������  �t$H��tj�|A�L$�@Q�@�С|A�L$�@V�@Q�D$H   �С|A�L$�@Q�@�D$L�����Ѓ���������H@��t�|AV�@Q�@�Ѓ��L$4d�    Y_^[��0� ��������VW��跻���t$�΍xH詻���H ���_^� �������������W��舻���x` u	� }  _� V���q����t$�ύp`�c����H ���^_� �������SVW���F����x` u� }  �$���2����p`�D$���P�������H ��Ћ��|A�\$�IS�I�у�;�@�|AS�@�@�Ѓ�;�+���ߺ���t$���t$�pDS�t$�Ⱥ���H ���_^[� _^�����[� W��診���xP u	�����_� V��葺���t$ ���t$ �pP�t$ �t$ �t$ �t$ �o����H ���^_� ���W���X����xT u	�����_� V���A����t$���t$�pT�/����H ���^_� ���W�������xX tV���
����t$�ύpX������H ���^_� ���$P�t$ �D$    �D$    �D$    �D$    �D$    �D$    ���  ����t,�$��t%�t$�|A�t$�@�t$�@X�t$Q�Ѓ����3��������������������������̡|AQ���   � ��Y���������������SUV��L$�F�.�V���    �;�~|�
W�@�+����ρ�  �yI���Au��u	�   +���|Ah�Hh�   ��    P��  U�ЋЃ���t�N�~_�^�^]��[� �F_�F^]��[� �^^][� �������������A    �A    �A    �����V��~ ��u�|A�v�@4� �Ѓ��F    �F    ^���������������̸   ����������̸   �����������3�� ������������ ������������̡|AV�@4��@$h�  �v���t$�|A�t$�@4�t$�@�t$�v�Ѓ�2�^� ����������������t$��t$�t$�t$�P� ��������3�� ����������̸   � ��������� �������������Q�|AU�@V�@ W�|$���3���=INIb�!  �  =SACbqt(=$'  t
=MicM�i  �E W���P$�   _��^]Y� �E �L$Q�L$Q�͉t$�t$�P��t�t$�|A�t$�@4�u�@�Ѓ��   _��^]Y� =ARDb�  �|AS�@j ���   j���Ћء|Aj �@j���   ���ЋL$���|Aj �@j���   �ЋL$��|Aj �@j���   ���t$�U PVWS���R[�   _��^]Y� �E ���P�   _��^]Y� =NIVb\tD=NPIbt-=ISIbuS�u ����  P���  P���V�   _��^]Y� �E W���P_^]Y� �E ���P�   _��^]Y� =cnyst	_��^]Y� �|Aj �@hIicM���   ���ЋU WP���R _^]Y� ������������j�h��d�    P��,V�8A3�P�D$4d�    ��~ ��   �|A�v�@4�@�Ѓ|$H t+�|AP�F�I0�p�Al�Ѓ��L$4d�    Y^��8� ���L$ hARDb�D$�D$    ��  �NP�D$P�D$P�D$H    �  �|A�L$���   Q� �Ѓ��L$ �D$<�������  �L$4d�    Y^��8� ����������̡|A�t$�@4�q�@l�Ѓ��   � ̡|A�q�@4�@�Ѓ�������������̡|A�q�@4�@�Ѓ�������������̡|A�q�@4�@�Ѓ�������������̡|A�q�@4�@|�Ѓ�������������̡|A�q�@4���   �Ѓ����������̡|A�t$�@4�q�@(�Ѓ�� �������t$�|A�t$�@4�t$�@,�q�Ѓ�� ���������������t$�|A�t$�@4�q�@0�Ѓ�� �̡|A�q�@4�@4��Y��������������̡|A�t$�@4�q���   �Ѓ�� ��̡|A�t$�@4�q�@ �Ѓ�� �����̡|A�t$�@4�q�@$�Ѓ�� �����̡|AV���   �t$�@WV���Ѓ����|AV���   u�@@�Ћ|AP�I4�w�A �Ѓ�_^� �@�Ѓ����|Au&���   V�@8�Ћ|AP�I4�w�A$�Ѓ�_^� �@h���0  h
  �Ѓ�_^� ����������������t$�|A�t$�@4�q�@D�Ѓ�� ���t$�|A�t$�@4�q�@H�Ѓ�� ���t$�|A�t$�@4�q�@L�Ѓ�� ���t$�|A�t$�@4�q�@P�Ѓ�� �̡|AS���   V�@W�|$W���Ѓ����|A���   �@��   �t$V�Ѓ����|AV���   u5�@@�Ћ|AW���   ���I@�ы|AV�I4P�s�AP�Ѓ�_^[� �@�Ѓ����|Au<���   V�@8�Ћ|AW���   ���I@�ы|AV�I4P�s�AH�Ѓ�_^[� �@h��0  h�  �Ѓ�_^[� W�Ѓ����|A��   ���   �t$�@V�Ѓ����|AV���   u5�@@�Ћ|AW���   ���I8�ы|AV�I4P�s�AL�Ѓ�_^[� �@�Ѓ����|Au<���   V�@8�Ћ|AW���   ���I8�ы|AV�I4P�s�AD�Ѓ�_^[� �@h4��0  h�  �Ѓ�_^[� �@hT��0  h�  �Ѓ�_^[� ����������t$�|A�t$�@0�t$���   �t$�q�Ѓ�� ������̡|A�t$�@0�q���   �Ѓ�� ����D$�|A���@0�$�t$���   �t$�q�Ѓ�� ��t$�|A�t$�@4�t$�@�t$�q�Ѓ�� �����������t$�|A�t$�@4�t$�@�t$�q�Ѓ�� �����������t$(�|A�t$(�@4�t$(�@T�t$(�t$(�t$(�t$(�t$(�t$(�t$(�q�Ѓ�,�( ���t$�|A�t$�@4�t$��  �t$�q�Ѓ�� ��������t$ �D$�t$ �|A�t$ �@4�t$ ��  ���D$�D$$�$�q�Ѓ�$�  ������������̡|Ah�����@4h�����@Th�����t$�t$h����h����h����h�����t$(�q�Ѓ�,� ����������̡|A�t$�@4�q�@8�Ѓ�� �����̡|A�t$�@4�q�@<�Ѓ�� �������t$�|A�t$�@4�q���   �Ѓ�� ��������������̡|A�q�@4�@@�Ѓ�������������̡|A�q�@4��  �Ѓ����������̡|A�D$�@4����  �$�q�Ѓ�� ����������t$�|A�t$�@4�t$�@X�t$�q�Ѓ�� ���������̡|A�q�@4�@`��Y��������������̡|A�q�@4�@d�Ѓ���������������t$�|A�t$�@4�t$��   �t$�q�Ѓ�� ��������t$�|A�t$�@4�t$�@\�t$�t$�t$�q�Ѓ�� ���t$�|A�t$�@4�q��  �Ѓ�� ����������������t$�|A�t$�@4�q�@h�Ѓ�� ���t$�|A�t$�@4�q��  �Ѓ�� ����������������t$�|A�t$�@4�q�@p�Ѓ�� ��j�h��d�    P��VW�8A3�P�D$ d�    ��hYALf�L$�[�  P�|A�w�B4�D$0    �@l�Ѓ��L$�D$(�����m�  �L$ d�    Y_^�� ������������UVW�|$���t�|A�L$�@j ���   j�Љ�t$��t�|A�L$�@j ���   j�Љ�|AV�@4W�u�@p�Ѓ�_^]� �������������t$�|A�t$�I�@0�t$���   �q�Ѓ�� ���������t$�|A�t$�@4�t$�@x�t$�q�Ѓ�� ���������̡|A�t$�@4�q�@t�Ѓ�� �������t$�|A�t$�@4�t$���   �t$�t$�q�Ѓ�� ����t$�|A�t$�@4�t$���   �t$�t$�q�Ѓ�� ��̃��|ASW�D$    �D$    �@�ًL$$���   �{j j�ЋL$$�D$�|Aj �@j���   �ЉD$�|A�L$�@0Q�@`�L$Q�w�С|A�s�@4�@�Ћ|Aj �I0�T$,R�T$4R�T$(R�T$4RP�C�p�Ah�Ѓ�,�|$( _[t.�|$$ t.�L$�T$;�~C�D$�;�}9�$�T$;�~.�D$��|$$ u�L$�T$;�~�D$�;�}�   ��� 3���� ����������������t$�D$�|A���@4�D$�D$���   �$�t$�q�Ѓ�� ������t$�|A�t$�@4�t$���   �q�Ѓ�� ����������̡|A�q�@4���   �Ѓ����������̡|A�q�@4��  �Ѓ�����������V��V���|AhP� �@0� �Ѓ��F�F    ��^�����V��N����t�|AQ�@0�@�Ѓ��F    ^������̸   ����������̸   ����������̸   � ��������3�� �����������3���������������� ����������������������������̡|AV�@W�|$�@ �����=NIVb��   ��   =TCAbttK=$'  t2=MicM��   �|Aj �@hIicM���   ���ЋWP���R_^� �W���P_�   ^� �|Aj �@hdiem���   ���ЋWP���R_^� =INIbuz�~ u���F   �P_^� �~ t�����P_^� =atni=t/=ckhct=ytsdu8����P_�F    3�^� ����P_^� ��  _3�^� =cnys����_3�^� �����V��N��u3�^� �|Aj �@0j ���   j j j �t$4j �t$(jQ���t$D�|A�t$D�@0�t$D���   �t$Dj �t$D�v�Ѓ�D^� ��������̋I��u3�á|AQ�@0�@�Ѓ�����̋I��u3�� �|AQ�@0�@�Ѓ�� j�h7�d�    P��V�8A3�P�D$d�    �D$    �q��u �D$,�    �p�L$d�    Y^�� � �D$0�H��|AQ�t$8�@0R���   �L$VQ�ЋЋt$@j �    �F    �|AR���   V�@�D$D   �Ћ|A�D$,���   P�	�D$,   �D$H �у�$�ƋL$d�    Y^�� � �������������̡|A�t$�@0�q���   �Ѓ�� ��̡|A�q�@0���   �Ѓ����������̡|Aj �@0j ���   j j j j j j j4�q�Ѓ�(�������̡|Aj �@0j ���   j j j j j j j;�q�Ѓ�(�������̡|A�t$�@0�q�@�Ѓ�� �����̋I��t(�|Aj �@0j ���   j j j j �t$j jQ�Ѓ�(� ���������������t$�|A�t$�@4�t$�@,�q�Ѓ�� ���������������t$�|A�t$�@4�q�@0�Ѓ�� �̡|A�q�@4�@4��Y���������������V�q��u3�^� �D$�H��|AQ�t$�@0R�@V�Ѓ�^� ��������������V�q��u3�^� �D$�H��|AQ�@0R���   V�Ѓ�^� ��������������̋D$3�h�����h  ���Pj BRj �t$ �t$ �   � ����j�hb�d�    P��$VW�8A3�P�D$0d�    ��htniv�L$ ���  �|A�t$D�@hulav�@4�L$$�D$@    �С|Ahgnlf�@htmrf�@4�L$$�С|A�t$H�@hinim�@4�L$$�С|A�t$L�@hixam�@4�L$$�С|A�t$P�@hpets�@4�L$$�С|A�t$T�@hsirt�@4�L$$�ЋL$X�t$\��  �u�����t.�|AQ�@h2nim�@4�L$$�С|AV�@h2xam�@4�L$$�ЍD$P�t$D�D$P������P�|A�D$<���   �@8�Ћ|A�����   �D$�	P�D$@ �у��L$�D$8�������  �ƋL$0d�    Y_^��0�  ��������������U����j�h��d�    P��pV�8A3�P�D$xd�    ��htlfv�L$4�V�  �|A�E�@���@,�$hulav�L$<Ǆ$�       �С|A�u,�@htmrf�@4�L$8�С|A�E�@���@,�$hinim�L$<�С|A�E�@���@,�$hixam�L$<�С|A�E$�@���@,�$hpets�L$<�С|A�uD�@hsirt�@4�L$8���U0W�f.џ��Dz�E8f.����D{A�|A���@�$�@,h2nim�L$<�С|A�E8�@���@,�$h2xam�L$<�С|A�u@�@hdauq�@4�L$8�ЍD$0P�u�D$$P������P�|AƄ$�   ���   �@8�Ћ|A�����   �D$ �	PƄ$�    �у��L$0Ǆ$�   ������  �ƋL$xd�    Y^��]�@ ����������t$(W�j ���D$�$�D$8htemf�� �D$�D$T�D$�D$L�D$�D$D�$�t$@�����( �������L$f.����%����D{�Y��^��T$f.����D{�Y��^��t$(W�j ���D$�$�D$8�Y�hrgdf�� �^��D$�D$D�L$�T$�$�t$@�����( ���t$(��W�j ���D$�$�D$8�^�htcpf�� �D$�D$T�^��D$�D$L�^��D$�D$D�$�t$@�����( ��U����j�h��d�    P��hSVW�8A3�P�D$xd�    �ًE��u)�|A�@���   �Ѕ�u�L$xd�    Y_^[��]� ����  htlfv�L$4��諷  �ufn�������YǄ$�       �D$�D$�$�< �F�\$$�D$�D$�$�< �D$$�\$�^D$�|A�$�@hulav�@,�L$<�С|Ahmrff�@htmrf�@4�L$8�Ћufn�������Y�D$$�D$$�$�+< �F�\$�D$$�D$$�$�< �D$�\$$�^D$$�|A�$�@hinim�@,�L$<�Ћufn�������Y�D$$�D$$�$��; �F�\$�D$$�D$$�$�; �\$$�D$�^D$$�|A�$�@hixam�@,�L$<�С|A���@���@,�$hpets�L$<�С|Aj �@hdauq�@4�L$8�С|AW�@hspff�@4�L$8�С|A�u �@hsirt�@4�L$8�ЍD$0P�u�D$$P������P�|AƄ$�   ���   �@8�Ћ|A�����   �D$ �	PƄ$�    �у��L$0Ǆ$�   ����赵  �ƋL$xd�    Y_^[��]� ��������������j�h��d�    P��$V�8A3�P�D$,d�    ��hCITb�L$��  �|A�t$@�@hCITb�@8�L$ �D$<    �С|A�t$D�@hsirt�@4�L$ �С|A�t$H�@hulav�@4�L$ �ЍD$P�t$@�D$P���q���P�|A�D$8���   �@8�Ћ|A�����   �D$�	P�D$< �у��L$�D$4����誴  �ƋL$,d�    Y^��0� �����V�q��u3�^� �D$�D$�H��|AQ�t$$�@0���@(�D$�D$(�$�t$$RV�Ѓ�$^� j�h�d�    P��V�8A3�P�D$d�    ��L$,�D$P����j �t$4��P�t$4�D$0    �b����|A���I�D$�IP�D$$�����у��ƋL$d�    Y^��� �������������V�q��u3�^� �D$�H��|AQ�@0�L$�@,QRV�ЋL$3҃�9T$^�� ��������������V�q��u3�^� �D$�H��|AQ�t$�@0R�@,V�Ѓ�^� ��������������V�q��u3�^� �D$�H��|AQ�t$�@0R�@0V�Ѓ�^� ��������������UVW���O����   �D$�l$�P�0�|AR�@0U�@0VQ�Ѓ���tb� t\�D$�H��|AQ�p0�EP�F0R�w�Ѓ���t6���t/�D$�H��|AQ�p0�EP�F0RW�Ѓ���t_^�   ]� _^3�]� �QV�q��u3�^Y� �D$W�H��|AQ�L$�D$    �@0Q�@8RV�Ћ�����t=�T$��t5�|A�t$�AR�@�Ћt$����t�|AV�@�@��V�&�������_^Y� �����������V�q��u3�^� �D$�H��|AQ�t$�@0�t$�@<RV�Ѓ�^� ���������̋D$��V���u�|A�@���   �Ѕ�u^��� W���O�  �v����t#�D$$�H��|AQ�@0�L$�@0QRV�Ѓ���fn�������Y��L$ �D$�D$�Y��$�>�  �~ �L$,_f��~@��f�A^��� ��������������j�h)�d�    P��V�8A3�P�D$d�    ��|A�L$�@Q�@�Ѓ��D$P�t$,���D$(    ��������t�L$,�D$P�ٙ���|A�D$�IP�I�D$$�����у��ƋL$d�    Y^��� ������V�q��u3�^� �D$�H��|AQ�@0j ���   j j j j j Rj1V�Ѓ�(^� ̡|AV�@j �t$���   ��L$��h���h  �j j jj P�t$$���%���^� ̡|AV�@j �t$���   ��L$���t$$���t$$j �t$(�t$(�t$(P�t$$�����^�  �������������U������<�|AV�@�����   W��$�u��M���\$8�E8j �u@�΃��D$�E0�$�u,�E$�� �D$�E�D$�E�D$�D$t�$�u�����^��]�< ���������������U������<�|AV�@�����   W��$�u��M���\$8j j ��W��D$�$�E$htemf�� ���D$�E�D$�E�D$�D$t�$�u�L���^��]�$ �����U������<�|AV�@�����   W��$�u��M���\$8�Uf.����%����D{�Y��^��Mf.����D{�Y��^�j j ��W��D$�$�E$�Y�hrgdf�� ���^��D$�D$t�T$�L$�$�u�x���^��]�$ �U������<�|AV�@�����   W��$�u��M���\$8��j W�j �����D$�$�E$�^�htcpf�� �D$�E�^��D$�E�^��D$�D$t�$�u�����^��]�$ ̃�0�|AV��W��D$���L$Q�t$H�D$�@�L$,���   Q�L$L���~ j �t$Tf�D$�t$T�~@�t$T�D$$P�t$P���t$Pf�D$8�����^��0� ���j�hT�d�    P�� V�8A3�P�D$(d�    ��|A�L$�@Q�@�Ѓ��L$<�D$P�t$D�D$ P�D$<    �v����t$D��j P�t$D�D$@�����|A���I�D$�IP�D$4 �ѡ|A�L$�@Q�@�D$8�����Ѓ��ƋL$(d�    Y^��,� ���j�h��d�    P��HV�8A3�P�D$Pd�    ��L$4�a����L$dP�t$l�D$ P�D$d    �J  �L$Q���D$\����j j P�t$l���D$h�`����|A���I�D$�IP�D$\�у��L$�D$X �����L$4�D$X�����Ԓ���ƋL$Pd�    Y^��T� ���������������U������x�U��V�uW���D$0���t.�|A���@W����   �$R�����\$0�D$0�D$0�|AW��L$8Q�u�D$@�D$H�D$P�@�L$p���   Q�����~ �wf�D$P�~@f�D$X�~@f�D$`��u
3�_^��]� �E�E�H��|AQ�u �@0���@(�D$�D$H�$�L$hQRV�Ѓ�$_^��]� ���V�q3���t,�D$�H��|AQ�@0�L$�@,QRV�Ћ�3���9D$���|AP�Q�t$�L$�R0�ҋ�^� �������������V�q��t#�D$�H��|AQ�@0�L$�@,QRV�Ѓ����|A�t$�A�t$�L$�@4�Ћ�^� ����̃�V�q��t#�D$�H��|AQ�@0�L$�@0QRV�Ѓ����|A�D$�A�L$�@,���$�t$ �Ћ�^��� ����̃�V�D$P�t$ W��t$ �D$���D$������|A���Q�L$ �R@�D$P�t$(�ҋ�^��� ������������̃�V��W�~W��D$�D$�D$����   �D$$�H��|AQ�@0�L$�@0QRW�Ѓ���t�~��tx�D$(�H��|AQ�@0�L$�@0QRW�Ѓ���tS�v��tL�D$,�H��|AQ�@0�L$�@0QRV�Ѓ���t'�|A�L$�@Q�t$8�L$8�@H��_�   ^��� _3�^��� �����������j�h��d�    P��V�8A3�P�D$d�    ��|A�L$�@Q�@�Ѓ��D$P�t$,���D$(    �����|A���Q�L$,�R8�D$P�t$4�ҡ|A�L$�@Q�@�D$$�����Ѓ��ƋL$d�    Y^��� ��������������j�h��d�    P��V�8A3�P�D$$d�    ��L$葌���D$P�t$8���D$4    �����|A���Q�L$8�R<�D$P�t$@�ҍL$�D$,�����;����ƋL$$d�    Y^��(� �����̃� V�qW��D$�D$�D$��t(�D$(�H��|AQ�@0�L$�@<Q�L$QRV�Ѓ����T$0���t�|A�A�L$�@HQ�L$0R�ЋT$4���t �|A�D$�@�L$,�@,���$R�Ћ�^�� � ����̋D$3҃8V�p�¸   h���h  ���E�3�����Rj @Pj V�t$$����^� �T$�t$3��:�t$��P�t$ �t$ �t$ �r�t$ ����� �T$�D$03��:��P�t$<���D$�D$@�$�t$<�D$8�� �D$�D$P�D$�D$H�D$�B�$�t$@�����8 ���̋D$3҃8�H��W�Rj ���D$�$�D$4htemf�� �D$�D$P�D$�D$H�D$�$�t$@�Q����  �������������̋D$�T$�h���%�3҃8��f.����D{�Y��^��L$f.����D{�Y��^�Rj ��W��D$�$�D$4�Y�hrgdf�� �^��D$�T$�L$�,$�t$@�����  ���������̋D$��3҃8W����PRj ���D$�$�D$4�^�htcpf�� �D$�D$P�^��D$�D$H�^��D$�$�t$@�����  ���������̋T$3��:��P�t$�B�t$�t$P�t$�t$�V���� ��̋D$�t$3҃8��RP�t$����� ���������������j�h�d�    P��$V�8A3�P�D$,d�    ��hgnrs�L$��  �D$@�D$4    �D$   �D$�|A�L$�@Q���   j�L$ �D$<�С|A�L$���   Q� �D$8 �ЋD$H���D$   �D$�|A�L$�@Q���   j�L$ �D$<�С|A�L$���   Q� �D$8 �Ѓ��D$P�t$@�D$P������P�|A�D$8���   �@8�Ћ|A�����   �D$�	P�D$< �у��L$�D$4�����P�  �ƋL$,d�    Y^��0� �����������W�y��u3�_� �D$�D$�H��|AV�p0�D$Q�t$(�����D$�D$,�$P�F(RW�Ѓ�$^_� ���������̡|Aj �@0j ���   j j j j j j j �q�Ѓ�(�������̋I��u3�� �|A�t$�@4�t$��  Q�Ѓ�� ����̋I��u3�� �|A�t$�@4�t$�@hQ�Ѓ�� �������̋I��u3�� �|A�t$�@4�t$�@pQ�Ѓ�� �������̋I��u3�� �|A�t$�@4�t$��  Q�Ѓ�� ������t$�|A�t$�@0�t$���   �t$�q�Ѓ�� ������̡|A�P0�D$�pj j j �t$�t$j �0���   j=�q�Ѓ�(� �����������̡|A�P0�D$�p�t$j j j��t$j �0���   j=�q�Ѓ�(� �����������̋D$�t$���PAEС|A�2�@0�t$�@@�q�Ѓ�� ��Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$jQ�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$jQ�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj �t$$�D$    �t$ �@0�t$ ���   �t$ �t$0�t$$jQ�ЋD$(��(Y� ��������������Q�I��u3�Y� �|A�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j*Q�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� ��Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� ��Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$j	Q�ЋD$(��(Y� ��Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$j
Q�ЋD$(��(Y� ��Q�I��u3�Y� �|A�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$j'Q�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$j,Q�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j:Q�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj j j �t$�D$    �t$ �@0j ���   j j)Q�ЋD$(��(Y� ������Q�I��u3�Y� �|A�$Rj j �t$�D$    �@0j �t$ ���   j j j)Q�ЋD$(��(Y� �����̋I��u3�� �|Aj �@0j ���   j �t$�t$�t$j �t$ jQ�Ѓ�(� ���Q�I��u3�Y� �|A�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j>Q�ЋD$(��(Y� Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� �̡|Aj �@0j ���   j �t$�t$�t$j �t$ j.�q�Ѓ�(� �������������V�q��u3�^� �D$�H��|AQ�@0j ���   j j j �t$ �t$(RjV�Ѓ�(^� �������������V�q��u3�^� �D$�H��|AQ�@0j ���   j j j j j RjV�Ѓ�(^� �V�q��u3�^� �D$�H��|AQ�t$�@0R�@\V�Ѓ�^� �������������̃�SVW�t$ �ٍL$�+�  �D$ P�D$P�L$�h�  ��tm�|$�L$ ��tJ�|AQ���   �@H�ЋS������tR�w�|Aj �A0j ���   j j �t$ V�7jR�Ѓ�(��t%�D$ P�D$P�L$���  ��u�_^�   [��� _^3�[��� ��������������Q�I��u3�Y� �|A�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� �̡|AV�@4W�|$� �w���ЋD$�G    �w�H��|AQ�t$�@0W���   R�v�Ѓ�3Ʌ����G_^��� �������̋I��u3�� �|Aj �@0j ���   j �t$�t$�t$j �t$ j/Q�Ѓ�(� ��̋T$��u3�� �r�B    �|A�t$�@0�q���   �Ѓ�� �����������̋I��u3�� �|Aj �@0j ���   j j j �t$j j jQ�Ѓ�(� ��������̡|Aj �@0j ���   j j j j j j j6�q�Ѓ�(�������̋I��u3�� �t$�|A�t$�@0�t$�@DQ�Ѓ�� ���̋I��u3��  �t$ �|A�t$ �@0�t$ ���   �t$ �t$ �t$ �t$ �t$ Q�Ѓ�$�  ������������̋I��u3�á|AQ�@0�@X�Ѓ�����̋I��u3�� �|A�t$�@0�t$�@LQ�Ѓ�� �������̋Q��u3�� �|A�H0�D$   �P�APR�Ѓ�� �����̋I��u3�� �|A�t$�@0Q�@P�Ѓ�� �����������̋I��u3�� �t$�|A�t$�@0�t$�@T�t$Q�Ѓ�� j�h+�d�    P��VW�8A3�P�D$ d�    ���L$��  �D$0�L$�P�0�|AR�@0Q���   j j j j j Vj8�w�D$P    �Ћ���(��t�L$4�D$P�2�  �L$�D$(������  �ƋL$ d�    Y_^�� � ����������̋D$V�P�0�|AR�t$�@0j ���   j j j j Vj9�q�Ѓ�(^� ���������̋D$V�P�0�|AR�t$�@0�t$�@h�t$�t$V�q�Ѓ�^� �������������UVW�|$���t�|A�L$�@j ���   j�Љ�t$��t�|A�L$�@j ���   j�Љ�|AV�@0W�u�@`�Ѓ�_^]� �������������t$�|A�t$�@0�t$���   �q�Ѓ�� ����������̋T$�|A�@0��t*���   R�q�Ћ|A�t$�ЋA0R���   �Ѓ�� �t$�@|�q�Ѓ�� �����t$�|A�t$�@0�t$�@p�t$�t$�q�Ѓ�� �������t$�|A�t$�@0�t$�@d�t$�t$�q�Ѓ�� �����̡|Aj �@0j �t$���   �t$ �t$ �t$j �t$ j3�q�Ѓ�(� ����������̋D$j ��|Aj �@0j ���   j j j j Rj�q�Ѓ�(� �D$j ��|Aj �@0j ���   j j jj Rj�q�Ѓ�(� �D$j ��|Aj �@0j ���   j j j j Rj�q�Ѓ�(� �D$V�P�0�|AR�@0j ���   j j j j j Vj"�q�Ѓ�(^� �����������̋D$V�P�0�|AR�@0j ���   j j j j j Vj5�q�Ѓ�(^� �����������̋D$V�P�0�|AR�@0j ���   j j j �t$ j Vj<�q�Ѓ�(^� ���������̡|AV�@0j ���   j j j j �t$ ��j �t$$j�v�С|A�t$8�@0�v�@t�Ѓ�0^� ��������̡|Aj �@0j ���   j j j j j j j�q�Ѓ�(�������̡|Aj �@0j ���   j j j j �t$j j�q�Ѓ�(� ��̡|Aj �@0j ���   j j j j j j j�q�Ѓ�(�������̡|Aj �@0j ���   j j j j j �t$ j�q�Ѓ�(� ��̡|Aj �@0j ���   j j j j �t$ �t$ j&�q�Ѓ�(� ̡|Aj �@0j ���   j j j j j j j(�q�Ѓ�(�������̡|Aj �@0j ���   j j j j j j j#�q�Ѓ�(�������̡|Aj �@0j ���   j j �t$�t$j �t$ j+�q�Ѓ�(� ��������������̡|Aj �@0j ���   j j j j j j j0�q�Ѓ�(�������̡|A�t$�@0�q���   �Ѓ�� ���j�hN�d�    P��V�8A3�P�D$d�    ���t$D�L$��  �|A�t$0�@h8kds�@4�L$�D$,    �С|A�L$DQ�L$Qj �t$L�D$T    �t$L�@0�t$L���   �t$L�t$Hj2�v�Ћt$l��(�L$�D$$����趌  �ƋL$d�    Y^�� � ̡|A�q�@0���   �Ѓ����������̋I��u3�� �|Aj �@0j ���   j j j j j �t$ j-Q�Ѓ�(� ��������̃��|AW�@j ���   ���L$(j�ЋL$$�D$�|Aj �@j���   �ЉD$�|A�L$�@0Q�@`�L$Q�w�С|A�T$�H0�D$,�pR�T$,R�T$$R�T$0R�0�Ah�w�Ѓ�(�|$( _t.�|$( t.�L$�T$;�~C�D$�;�}9�$�T$;�~.�D$��|$( u�L$�T$;�~�D$�;�}�   ��� 3���� ��SV�t$W��u�q�|A�\$�@j ���   hdiuM���Ћ���tH;>u_^3�[� �|Aj �@hIicM���   ����;�u�|Aj �@h1icM���   ���Шu��>_^�   [� ������������j�hq�d�    P��V�8A3�P�D$d�    �|A�t$,�@hfnic�@T���ЋЅ�t�|Aj
�A�ʋ��   �Ѕ���   hfnic�D$P����(  �t$0P���D$(    �L�  �L$�D$$�����+�  �|A�΋@�@ �Ѓ��t�|A�΋@�@ �Ѕ�u�|Ahfnic�@�΋@$�С|A�t$4�@j
�@8���ЋL$d�    Y^�� ����������̡|A�q�@0���   �Ѓ�����������j�h��d�    P��$V�8A3�P�D$,d�    ��hmnrs�L$�,�  �|A�t$@�@j�@4�L$ �D$<    �ЍD$P�t$@�D$P������P�|A�D$8���   �@8�Ћ|A�����   �D$�	P�D$< �у��L$�D$4������  �ƋL$,d�    Y^��0� ������������j�h��d�    P��$V�8A3�P�D$,d�    ��|$@ �SSSS�DSSSE�P�L$�N�  �|A�L$�@�D$4    �@ �Ћ|Aj�QP�B4�L$ �ЍD$P�t$@�D$P�������P�|A�D$8���   �@8�Ћ|A�����   �D$�	P�D$< �у��L$�D$4������  �ƋL$,d�    Y^��0� ���������������V��V���|AhP� �@0� �Ѓ��F�F    ���F   �F    ��^�V��N����t�|AQ�@0�@�Ѓ��F    ^�������V��N�F    ��tk�|Aj �@0j ���   j j j j j j jQ�С|A�t$<�H0�t$<3�9D$H�t$<���t$<j ��
P�v���   �Ѓ�D��t�~ t	�   ^� 3�^� �������������̋D$�A�I��u3�� �|AQ�@0�@�Ѓ�� ��������̡|AS�@�\$�@ V�����=ckhc��   tz=cksata=TCAb��   �|AW�@j ���   hdiem���Ћ��SW���F   �R�~ ��t��t��u3�������P�L���_^��[� �~ tg����P^[� �~ tU�|Aj �@0j ���   j j j j j j j �v�Ѓ�(��t)�F    ^�   [� =atnit�t$��S�\���^[� ^3�[� U��} ��   S�\$V�t$W�|$$��wy�$�� 9t$��   �f9t$��   �Z9t$��   �N9t$��   �B�D$;�~:;���   �0�D$;�|(;�~~�"�D$;�|;�|p��D$;�~;�~b�9t$uZ�|Aj �@0j ���   j j j j j �t$0j�u��fn������(j���D$fn�����$S趏  ���E    _^[]� �H� T� `� l� x� �� �� �� �� W��� �\  V�t$����   �$��� �D$f/D$�4  ��   �D$f/D$�  ��   �L$f/L$�  �   �L$f/L$��   �   �T$f/T$��   �D$$f/���   �n�T$f/T$r`�D$$f/���   �N�T$f/T$r@�D$$f/���   �.�T$f/T$v �D$$f/�sl��D$f.D$���DzX�|Aj �@0j ���   j j j j j �t$(j�w���D$L��(�t$,���D$�D$0�$V�"�  ���G    ^_�$ �I b� y� �� �� �� �� � "� >� �������������D$j���D$�D$0�D$�D$(�$�t$$�t$$�+����  ���������D$j���D$�D$0�D$�D$(�$�t$$�t$$������  ���������D$j���D$�D$0�D$�D$(�$�t$$�t$$�����  ��������V��V���|AhP� �@0� �Ѓ��F�F    �$�F   ��^��������V��N����t�|AQ�@0�@�Ѓ��F    ^������̡|AV�@��L$�@ ��=cksat]=ckhct�t$���t$�/���^� j j j j j j �F   �|Aj �@0j ���   j �v�Ѓ�(��t!�F    �   ^� �~ t����P^� 3�^� �j�h��d�    PQV�8A3�P�D$d�    ��t$���|AV�@0hP� � �Ѓ��F�F    �F   �D$ �L$�L�F�|Aj �@hmyal���   �D$    �ЉF��t��t�F    �|A�L$�@j
���   hhfed�ЉF�ƋL$d�    Y^��� ����̡|AV�@��L$�@ ��=ytsdt�t$���t$�v���^� �|A�v�@0���   �Ћ�����P�   ^� ������������3���������������3�������������������������������3���������������3���������������3���������������3�� �����������Q�L$�$    �o  �D$Y� ������̋A��uË ���������������������V���PD��t�D$9Ft
�F����PH^� ������������̋A�������������j0�t$���  ����j0�t$�5Q����P�܃  �����������j�h�d�    P���8A3�P�D$d�    �t$(�D$�t$(P�Q��j0P�D$0    苃  �|A�L$�@Q�@�D$4�����Ѓ��L$d�    Y�����������������j�h0�d�    P���8A3�P�D$d�    �t$,�D$�t$,�t$,P�gR��j0P�D$4    ��  �|A�L$�@Q�@�D$8�����Ѓ��L$d�    Y�������������j$�t$�ł  3Ƀ���������������j$�t$��O����P蜂  3Ƀ����������������������j�hS�d�    P��S�8A3�P�D$d�    �t$,�D$�t$,P��O��j$P�D$4    �:�  �|A3ۋI���I�D$P���D$8�����у��ËL$d�    Y[����j�hv�d�    P��S�8A3�P�D$d�    �t$0�D$�t$0�t$0P�Q��j$P�D$8    趁  �|A3ۋI���I�D$ P���D$<�����у��ËL$d�    Y[���������������̡|A�t$�@�t$���   j �Ѓ�����t$�|A�t$�@�t$���   j �Ѓ���������������̡|A�@���  ��|A�@0���   ��j�h��d�    P��VW�8A3�P�D$ d�    �t$8�D$    �|A�t$8�@0�L$���   Q�Ћ��|A�|$<�IW�I�D$8   �ѡ|AW�@V�@�Ћ|A�D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� ����j�h��d�    P��(SUVW�8A3�P�D$<d�    �D$    �|A�|$L�@W�@�D$H    �Ѓ��|A�L$P�@3ۋ��   SS�D$L    �D$    �ЋL$P�D$�|AS�@j���   �Ћ����&  3���I ��~|�|A�L$�@Q�@�С|Aj �@j��@�L$(hxQ�Ѓ��|A�ϋ@�D$D   �@<�Ћȡ|Aj��@j��@L�T$$RQ���С|A�L$�@Q�@�D$H �Ѓ�V�t$�D$4P�!�������|A�ϋ@�D$D   �@<�Ћȡ|Aj��@j��@LVQ���С|A�L$,�@Q�@�D$H �С|A�L$T�@�����   j ��
UC�ЉD$�|Aj �P�M���   Q�L$X�ҋ���������ǋL$<d�    Y_^][��4�����������̡|A�@0���   ��|A�@0���   ��|A�@0���   ����W��JR��A(�P$j j h������  �������������̸|�����������j�hA�d�    P��8SVW�8A3�P�D$Hd�    ����L$Q���P(���W�D$P    ��t&�|Aj �A0j ���   j j j j Vj jR�Ѓ�(�|A�L$�@Q�@�D$T�����С|A�L$�@Q�@�Ѓ��O�D$P   ��t'�|Aj �@0j ���   j �T$ Rj jj?j Q�Ѓ�$�|A�L$�@Q�@�D$T�����С|A�L$�@Q�@�Ѓ��O�D$P   ��u3��>�|A�T$Rj j j h  
 j�T$,R�D$,    �@0h�  ���   jQ�ЋD$8��(���|A�L$�@Q�@���D$T�����Ѓ���t3��L$Hd�    Y_^[��Dá|A�L$�@Q�@�Ѓ��O�D$P   ��t'�|Aj �@0j ���   j �T$ Rj j j8j Q�Ѓ�$�|A�L$�@Q�@�D$T�����ЋO����t�|Aj�@0Q�@P�Ѓ��L$4�v  ���|A�D$$�IP�I�D$T   �у�Vh   h  K j;�D$4Ph	��h�  ���D$l�R����|A�L$$�@Q�@�D$T�Ѓ��L$4�D$P�����v  �O��t�|AQ�@0�@X�Ѓ��O��t�|AQ�@0�@X�Ѓ��O��t&�|Aj �@0j ���   j j j jj j jQ�Ѓ�(j�$�`z  ���   �L$Hd�    Y_^[��D������j�hd�d�    P��VW�8A3�P�D$$d�    ��j�N��  �F4    �F8    �F<    W��F(�|Ah�   �@0�v�@�С|A�L$�@Q�@�С|Aj �@j��@�L$(h�Q�Ѓ�j j �D$P�D$P���D$<    �D$�  �D$     谿���|A�L$�@Q�@�D$0�����Ѓ��Nj j��  �L$$d�    Y_^��$������j�h��d�    P��\VW�8A3�P�D$hd�    ��|A�L$�@Q�@�С|Aj �@j��@�L$ h�Q���F(�Y�Ǆ$�       �D$ �  �D$$    �,�P�D$LP��8���L$0QP�D$HPƄ$�   �  ��(j j P�D$P��Ƅ$�   豾���|A�L$$�@Q�@�D$t�С|A�L$8�@Q�@�D$x �С|A�L$�@Q�@�D$|�����Ѓ��L$Thtats�s  �|Aj�@j�@0�L$\�D$x   �С|A�F(�@�@,���L$\�$j�ЍD$TP�D$P�D$LP���D$�  �D$    �����|A�L$D���   Q� �Ѓ��~4 t_�|A�N0�@P�@h�ЋF4��t�v8�Ѓ��F<�F8    �F4    ��|Ah��@h�  ��0  �Ѓ��|A�N0�@P�@l�ЍL$T�D$p������r  �L$hd�    Y_^��h� ����j�h��d�    P��@VW�8A3�P�D$Ld�    ��|A�|$\�@�ϋ@ ��=MicM��   =ckhctg=fnic�9  j�L$<�>r  �L$`P�D$X    �|r  �L$8�D$T�����[r  �|A�L$`�@j�@4j�и   �L$Ld�    Y_^��L� ����P����؋L$Ld�    Y_^��L� �|Aj �@hIicM���   ����=�����   htats�L$(�q  �|Aj �@j�@0�L$,�D$\   �ЍD$$P�D$P�D$P���D$�  �D$    �����|A�L$���   Q� �Ѓ��L$$�D$T�����oq  �N�F   ��t�|AQ�@0�@�Ѓ��t$`��W�����L$Ld�    Y_^��L� �l$V��t3�^� j�N�6�  j�Ou  �N���F    ��t�|AQ�@0�@�Ѓ��   ^� ����j�����  j�u  ��3������������D$�A(� �̍A�������������VW��~4 tC��    �|Ah��@h~  ��0  ��j
�  �|A�v �@P�@�Ѓ���uM9F4uá|A�N0�@P�@h�Ѓ~4 t9�|Ah��@h�  ��0  �С|A���@P�N0�@l���o���_3�^� �D$�F8�D$�F4�|AS�@P�N0�@l�Ѓ~4 t#j
�  �|A�v �@P�@�Ѓ���u89F4uݡ|A�N0�@P�@h�Ћ~<�F<    �|A�N0�RP�Rl��[��_^� [_3�^� �j�h��d�    P��V�8A3�P�D$d�    �L$��n  �L$0�|A�D$$    ��t"�@4Q�@�Ѓ���t'��L$Q�t$8���R(�'�@0�t$,�@�Ћȃ���u3��?��T$R�t$8�P ��|A�L$�@�@ �Ѓ��t�|A�L$�@0Q�t$0�@x�Ѓ��L$�D$$�����n  �ƋL$d�    Y^�� á|AV�@j �t$���   ��L$�Ћ���u�    �F^� ��u9Ft�   ^� ������������V�t$W��;t$u�|A�L$�@j ���   htsem�Ѕ�u`�|A�L$�@j ���   hrdem�Ѕ�uA�D$�D$�H��t2�|Aj �@0�T$�@,RVQ�Ѓ���t�t$���M
  _�   ^� _3�^� ������������j�h �d�    P��0VW�8A3�P�D$<d�    ���|A�L$�@Q�@�С|A�L$ �@Q�@�D$L    �Ѓ��L$L�D$P�t$T�D$4P�D$P��P���Ћ|A�D$D�A�L$�@QR�С|A�L$4�@Q�@�D$P�С|A�L$(�@Q�@�D$T �С|A��@V�@�С|A�L$ �@V�@Q�Ѓ����
  �|A�L$�@Q�@�D$H�����Ѓ��L$<d�    Y_^��<� �������j�hC�d�    P��SV�8A3�P�D$$d�    �ًt$<;t$@��   �|A�L$8�@j ���   htsem�Ѕ���   �|A�L$8�@j ���   hrdem�Ѕ���   �|A�L$�@Q�@�Ѓ��L$4�D$P�D$P�D$4    �t$�D$    虹����u3��5�|A���@��@V�С|A�L$(�@V�@Q�Ѓ����a	  �   �|A�D$�IP�I�D$0�����у��ƋL$$d�    Y^[��$� 3��L$$d�    Y^[��$� �̡|AV�@j �t$���   ��L$�Ћ���u�    �F^� ��u9Ft�   ^� �����������̃�V�t$W��;t$ uy�|A�L$�@j ���   htsem�Ѕ�uZ�|A�L$�@j ���   hrdem�Ѕ�u;�L$�D$�D$�D$P�D$P�t$������t�t$���  _�   ^��� _3�^��� �����������̃��|AV�@�����   W��$�t$��L$���\$����u�D$�    �F^��� ��u�Ff.D$���D{�   ^��� �̃�SV�t$��;t$ ��   �|A�L$�@j ���   htsem�Ѕ�ur�|A�L$�@j ���   hrdem�Ѕ�uS�D$W��H�D$��t?�|Aj �@0�T$�@0RVQ�Ѓ���t"�D$�����$�  ^�   [��� ^3�[��� ��0�|AV��W��L$Q�t$@�D$�D$�D$�@�L$$���   Q�L$D���~�~P�~H����uf�^f�V�    f�N^��0� ��u3�Ff.ß��Dz�Ff.��Dz�Ff.����D{�   ^��0� ���̃�4�D$@S�\$HV�t$TW�|$T�L$;�t;�t;���   �|A�L$H�@j ���   htsem�Ѕ���   �|A�L$H�@j ���   hrdem�Ѕ���   �L$D�D$�D$�D$$�D$(P�D$P�D$ PW��D$,P�D$8�D$@�D$H�t$ �|$(�\$0�������t<�~D$(�L$����f� �~D$Hf�@�~D$Pf�@�  �   _^[��4� _^3�[��4� ����������̃�0�|AV��W��D$���L$Q�t$@�D$�@�L$,���   Q�L$D���~ �~H�f�D$f�L$���uf�F�    f�N^��0� ��u�D$P�FP�  ����t�   ^��0� �������̃�SV�t$0��;t$4��   �|A�L$(�@j ���   htsem�Ѕ���   �|A�L$(�@j ���   hrdem�Ѕ�uh�L$$�D$�D$P�t$0W��D$���D$P�D$$�t$������t.�~D$���ċ�f� �~D$(f�@�  �   ^[��� ^3�[��� �������j�hs�d�    P��V�8A3�P�D$d�    ��t$�V�    �B    �D$$    ������D$    �D$    �|Aj ���   �L$�@QR�D$0�С|A�L$���   Q� �D$4 �Ѓ��ƋL$d�    Y^�� ������������̃�V�t$W�|$ �f.���Dz�Ff.G���D{a�G�Y����D$�D$�$��  �F�\$�Y�D$�D$�$���  �D$�\$��f.D$���D{_�   ^���_3�^���������������j�h��d�    PQV�8A3�P�D$d�    �D$    �|A�t$�@V�@�D$    �С|AV�@�t$(�@�Ѓ��|A�΋@�D$    �@<�D$   �Ћ|Aj��Qj��t$,�RLP���ҋƋL$d�    Y^���������������V��~ ��u�|A�v�@4� �Ѓ��D$�F    �F    t	V�42������^� �����������V��N����t�|AQ�@0�@�Ѓ��D$�F    t	V��1������^� �̋���u�D$�    �A� ��u�A;D$t�   � ��̋���u�D$�    �A� ��u�Af.D$���D{�   � ������̋���u*�~D$f�A�~D$f�A�~D$�    f�A� ��u9�Af.D$���Dz"�Af.D$���Dz�Af.D$���D{�   � ���������������V�����u �~D$f�F�~D$�    f�F^� ��u�D$P�FP���������t�   ^� ���j�h��d�    PV�8A3�P�D$d�    ���D$    ���u!�    �|A�N�@Q�@�L$Q�Ѓ��#��u�|A�T$�@�N�@xR�Ѕ�t�   �|A�L$�@Q�@�D$�����Ѓ��L$d�    Y^��� ����������j�h!�d�    P���8A3�P�D$d�    �t$0�D$    �|A�T$�@R�@P�ЋL$,P�D$(   �a  �L$�D$   �D$$ �'a  �D$,�L$d�    Y��$� �j�ha�d�    P�� �8A3�P�D$$d�    �t$<�D$    �|A�t$<�@�T$���   R�ЋL$4P�D$0   �VH���L$�D$   �D$, ��H���D$4�L$$d�    Y��,� ���������̡|A�D$�@H���@�$Q�Ѓ�� �������������̡|Aj �@HQ���   �Ѓ����������̡|A�t$�@Hj ���   Q�Ѓ�� ��̡|Aj�@HQ���   �Ѓ����������̡|A�t$�@Hj���   Q�Ѓ�� ��̡|Aj�@HQ���   �Ѓ���������̡|A�t$�@Hj���   Q�Ѓ�� ��̡|AQ�@H���  �Ѓ������������̡|A�t$�@HQ���  �Ѓ�� ����̡|A�t$�@HQ���  �Ѓ�� ����̡|A�t$�@HQ���  �Ѓ�� ����̡|A�t$�@H�t$��  Q�Ѓ�� ̡|A�t$�@H�t$��  Q�Ѓ�� ̡|AQ�@H���   �Ѓ�������������VW�t$���Ӭ  ������t�|A�t$�AHV���   W�Ѓ���_^� ���������VW�t$���t$�O�  ������t�|A�t$�AHV���   W�Ѓ���_^� ����̡|A�t$�@H�t$���   Q�Ѓ�� ̡|A�t$�@H�t$���   Q�Ѓ�� ̡|A�t$�@HQ���   �Ѓ�� ����̡|AQ�@H���  �Ѓ��������������t$�|A�t$�@H�t$���  �t$�t$Q�Ѓ�� �����j�h��d�    P��VW�8A3�P�D$ d�    ���|Aj �@Hh�  ���   W�Ѓ��|$0 ��   h�  �Y�  ��������   �|Aj �IHV���   W�у��L$�\  �|A�t$4�@h�  �@0�L$�D$0    �С|A�D$8�@���@,�$h�  �L$�С|Aj �@@�L$�@(QV�Ѓ��L$�D$(�����\  �   �L$ d�    Y_^�� � 3��L$ d�    Y_^�� � ������������̡|AQ�@H���   ��Y�������������̡|A�t$�@HQ���  �Ѓ�� ����̡|A�t$�@HQ���  �Ѓ�� ����̡|AQ�@H��4  �Ѓ������������̡|A�@H� �����̡|AV�@@�t$�@�6�Ѓ��    ^��S�\$U�l$V�}  W��u3�|AS�@HW���   �Ѓ���u�|Aj�@HW���   �Ѓ���t�   �t$�E ����   �|AW�@H���   �Ѓ��|$( u!�t$$�|AU�t$$�@HV���  SW�Ѓ��D��t@��I �t$$�|AU�t$$�@HV���  SW�С|A�����   �΋@(�Ћ���uɋt$�}  u�|AW�@H���   �Ѓ���t3���   �E ���|AW�@Hu$���   �С|AS�@HW���   �Ѓ�_^][� ���   �С|A���|$( �@Hu!�t$$���  j �t$$VSW�Ѓ���_^][� � h  �Ћ����u_^][� �|A�΋��   �@x�Ћ|AP���   �͋B|�Ѕ�tP�t$$�|Aj �t$$�@HV���  SW�Ћȃ���t�|AU���   �@H�С|A�΋��   �@(�Ћ���u�_^��][� ����t$�|A�t$�@H�t$���  �t$�t$Q�Ѓ�� ����̡|AQ�@H���   ��Y�������������̡|AQ�@H���   �Ѓ������������̡|A�t$�@H�t$���   Q�Ѓ�� ̡|AQ�@H���   ��Y�������������̡|AQ�@H��t  ��Y�������������̡|AQ�@H��P  �Ѓ������������̡|AQ�@H��T  �Ѓ������������̡|AQ�@H��X  �Ѓ������������̡|A���@HQ��\  �L$Q�ЋL$$�~ f��~@f�A�~@f�A���� � ��������������̡|AQ�@H��`  �Ѓ������������̡|A�t$�@HQ��d  �Ѓ�� ����̡|A�D$�@H����h  �$Q�Ѓ�� ����������̡|A�D$�@H����t  �$Q�Ѓ�� ����������̡|A�D$�@H����l  �$Q�Ѓ�� ����������̡|A�t$�@HQ��p  �Ѓ�� ������t$�|A�t$�@H�t$���  �t$Q�Ѓ�� ����������t$�|A�t$�@H�t$���  �t$�t$�t$Q�Ѓ�� ̡|Ah�  �@H� �Ѓ������������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@H���   �Ѓ������������̡|AQ�@H���   �Ѓ������������̡|A�t$�@HQ���   �Ѓ�� ����̡|A�t$�@HQ���   �Ѓ�� ����̡|A�t$�@H�t$���  Q�Ѓ�� ̡|A�t$�@H�t$��   Q�Ѓ�� ��t$�|A�D$�@H�����  �$Q�Ѓ�� ������̡|AV�@Hh  � �Ћ�������   �t$h�  �S�  �Ѓ���t^�|Aj �AHR���   V���t$h(  �'�  �Ѓ���t2�|Aj �AHR���   V�С|A�����   j �@j���Ћ�^á|AV�@@�@�Ѓ�3�^�������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@H��  �Ѓ������������̡|AQ�@H��  �Ѓ������������̡|AQ�@H���  �Ѓ������������̡|AQ�@H���  �Ѓ������������̡|AQ�@H���  �Ѓ������������̡|A�t$�@H�t$��  Q�Ѓ�� ��t$�|A�t$�@H�t$��   Q�Ѓ�� ��������������t$�|A�t$�@H�t$��|  �t$Q�Ѓ�� ��������̋D$V���u�|A�@H���  �'��u�|A�@H���  ���u(�|A�@H���  V�Ѓ���tP�t$���   ^� 3�^� ������������̃�SW���$�  �؅��  �|$$ �  �|AV�AHj ��p  h�  W�Ћ|A���IHh�  ���   W�t$0�������D$��u^_��[��� �|$(U3�ωl$�m�  ����   ��I �D$P�D$ P�t$ ��U�*�  ��tf�t$;t$\�l$ ������u����ɋD�;D�t.�|A�Hl����P�D$,�p�A�ЋD������tP����  F;t$~��l$�|$,E�ωl$�ԧ  ;��l���]^_��[��� _3�[��� �����̃��|AU�@Hj ��p  ��h�  U�l$�Ѓ��D$��u]��� �D$W��u�|A�@H���  �+��u�|A�@H���  ����Z  �|A�@H���  U�Ћ������<  S��蟧  �|Ah�  �@H3ۋ��   U�\$(�Ѓ�����   �l$V�s���|A�L$�@lS�q�@�Ћ؃�����   �|A�s�I\�t$$�I,�у���t�F�P���Ħ  �|A�s�@\�t$$�@,�Ѓ���t�F�P��螦  �E ;Et#�|A�s�@\�t$$�@,�Ѓ���tV���s�  �|A�s�@\�t$$�@,�Ѓ���t�FP���M�  �|A�\$$�@Hh�  �t$���   C�\$,�����Ѓ�;�����^[_�   ]��� _3�]��� ̡|AQ�@H���  �Ѓ������������̡|A�t$�@H�t$���  Q�Ѓ�� ��t$�|A�t$�@H�t$���  Q�Ѓ�� ������������̡|AQ�@H���  �Ѓ������������̡|AQ�@H���  �Ѓ������������̡|A�t$�@HQ��  �Ѓ�� ����̡|A�t$�@HQ��  �Ѓ�� ����̡|AQ�@H��  �Ѓ������������̡|A�t$�@HQ��  �Ѓ�� ����̡|AQ�@H��T  �Ѓ������������̡|A�t$�@H�t$��  Q�Ѓ�� ̡|A�t$�@HQ��8  �Ѓ�� ����̡|A�t$�@HQ��<  �Ѓ�� ������t$�|A�t$�@H�t$��@  Q�Ѓ�� ������������̡|A�t$�@HQ���  �Ѓ�� ����̡|A�t$�@HQ��H  �Ѓ�� ����̡|AQ�@H��L  ��Y�������������̡|AV�@Hh�  � �Ћ�����u^á|A�t$�@H�t$��  V�Ѓ���u�|AV�@@�@�Ѓ�3���^������������̡|AV�@@�t$�@�6�Ѓ��    ^���t$�|A�t$�@H�t$��   Q�Ѓ�� ������������̡|A�D$�@H����$  �$Q�Ѓ�� ����������̡|AQ�@H��(  �Ѓ������������̡|A�t$�@H�t$��,  Q�Ѓ�� ̡|A�@H��  ��|A�@H��  ��|AV�@@��@,WV�Ћ|A���ȋBj ���   h�  �Ћ|Ah�  �IHV���   ���у���
��t_3�^Ë�_^�̡|AQ�@@�@,�Ћ|A���ЋAj ���   h�  ������̡|A�D$�@H����  �t$,�t$,���$Q�L$Q�ЋL$4�~ f��~@f�A�~@f�A����0� ��������̡|A�D$�@H����  �t$,�t$,���$Q�L$Q�ЋL$4�~ f��~@f�A�~@f�A����0� ��������̡|AQ�@H���  �Ѓ������������̡|A�t$�@H�t$��8  Q�Ѓ�� ��t$�|A�D$�@H����0  �$�t$Q�Ѓ�� ��̡|A�@H�@����̡|AV�@@�t$�@�6�Ѓ��    ^���t$�D$�t$�|A���@H�$�t$���   �t$�t$�Ѓ�������������t$�D$�|A���@H�$�t$���   �t$�t$�Ѓ�����������������    ���������̡|Aj�@H�1��|  �Ѓ���������̡|AV�@H�t$��x  ����3Ƀ������^��� ������̡|Aj �@H�1��|  �Ѓ����������fnD$�L$����YD$�X��,�;�}���;D$OD$���������������̃�D�|AS�@HV���   W�|$Th�  W�Ћ|A3��IHV���   ��h�  W�\$L�у��D$L�t$�t$�t$��u
_^�C[��Dá|AU���   �ϋ@��=�  �|A�4  �@Hj ���   h:  W�Ћ|Ah�  �IHW���   �D$4�ы|A3�IHU���   h�  W�D$L�ы|A�؋IHW��  �\$H�ы|AW�IH�D$h���  �у�(3��D$D9t$,~z�K�ًD$@��tPj�W��謹  ���tA�L$D�@�|� ���L$L~�� ��%�������;�u&�(�  �L$L;�O���  ���;Cu�����G��;|$,|��\$$�D$ �|$X����   j W����  ����  �L$ 辛  ��tc�L$ �!�  �L$<;�uR�|A�I�@h����  ��h�  Q�L$X�Ѓ��D$H�D$����  �L$ �h�  �t$LP�t$P�T�  ���D$<h �@�|A���@h�  ���  Q�L$X�Ѓ��D$���<  �t$L�t$TP��  ����~-�|AhH�@h�  ���   ��U�Ѓ��D$����  �|Aj��@HV��  W�Ѓ�����  �l$ ��t!jW����  ����  ��轚  ���D$0�3��t$0�|Aj �@Hh�  ���   W�Ћ�3�3���T$ �l$(�D$89D$,�n  �{�|$<��L$@���z  j�P蜷  ����e  �L$D�@�|� �4��t$L~�� ��%�������9D$8��  ���ܳ  3�3��D$P�D$4    9^��   �l$$��������Шtm�D$������������������D$���T��N�D$�L��D$�J�L��N�D$�L���D$�J�L��N�D$�t$L�L���D$�J�L��C;^�y����l$(���<  �Ǚ+�����~�L$QPQ�L$�P  �\$ �L$0�m    �3��Ë�+ÉD$H�T$L��;D$P�  �D$����t3�D$�l$H�[�~�f�*�~D�f�D*�~D��ŋl$(f�D�D$�[�~�f��~D�f�B�~D�f�B;�}_�D$9�uR�L�����������w4�$��L$$��,��"�L$$��l���L$$��l��
�L$$��l���;�|��T$L�D$4�L$0E��@�l$(�T$L�D$4;�����;D$P�-  �|$<�T$ �D$8�t$0@���D$8�|$<;D$,������D$P�����D$ P�������  �T$ ��L$3�;G�Å���   �m    ōƋG��@�~�f��~D�f�B�~D�f�B�G��@�D$�~�f�B�~D�f�B �~D�f�B(��T$ �@�D$�~ȍȍm    �f�D�0�~Af�D�8�~Af�D�@��t7�G�@�D$�~ȍȍm    �f�D�H�~Af�D�P�~Af�D�X�G��@�D$�~ȍȍm    �f���~Af�D��~Af�D��G��o��@�D$E�~ȍȍm    �f���~Af�D��~Af�D���o��@�D$E�~ȍȍm    �f���~Af�D��~Af�D��/E�l$(��tC�G�@�D$�~ȍȍm    �f���~Af�D��~Af�D��oE�l$(�������G������D$P����D$ P����D$P�����3�]_^[��DË��   �ϋ@��=  ��  �|Aj �@Hh(  ���   W�Ћ|Ah(  �IHW���   ���ы��3ɉl$H��~�˅�t�|� �4Vu���A;�|�D$<hp�@�|A���@hY  ���  Q�L$X�Ѓ��D$����   �t$L�t$TP���  �|Ah��@��    ���  h^  Q�Ѓ��D$(��tL��    QSP��  �|A�ƋIH���   +���PVW�D$X�у���u!�D$P�u���D$,P�k����]_^3�[��Dá|Aj �@Hh�  ���   W�Ћ|Aj �IHh(  ���   W�D$h��3�3ۃ���3҉L$D�t$L�\$<���  �|$(��    �߅���   3��~y�L$P�R�4v�]�����D$C�~f��~Df�A�~Df�A�D$���~Df�A�~D f�A �~D(�D$<f�A(�|$(E�I0�v;�|��t$L�؃|� tg�|$P�.�@�D$�~ȍȍRBf���~Af�D��~Af�D��D$�v�~ȍȍRBf���~Af�D��~Af�D��|$(4ߋl$H�t$LC�\$<;�������L$D�T$@3���~��D�    ��   @;�|�D$(P�������D$P������   ]_^[��DÐ]ht������t$�D$�|A���@H�$�t$���  �t$�Ѓ���̡|A�@H���  ��|A�@H���  ���t$,�D$(�|A���@H�$�t$,���  �t$,�t$,�t$,�t$,�t$,�t$,�t$,�Ѓ�,����������̡|A�@H���  ��|A�@H���  ���t$,�D$�t$,�|A�t$,�@H�t$,��P  �t$,���D$�D$0�$�t$,�t$,�Ѓ�,����������A    ����q���|A�@l�@��Y��������̡|AV�@l��@�v�ЋL$����u	�   ^� �t$�|A�t$�@lQ�t$� ��3Ƀ������F^��� ������������̋I��u3�á|AQ�@l�@�Ѓ�����̃��|A�$�@lR�@�T$R�t$�t$�q�ЋL$�T$(��;�u	�$��� ���9$D���� ����̡|A�@H���   ��|A�@H���  �����|A�L$�@�����   W��$�t$���$�D$�$f/�w�D$f/�w(��|A�L$�@���@,�$�t$�Ѓ�������̃�0�|AW��$Q�t$<�D$�D$�D$�@�L$ ���   Q�L$@���~X�D$<f/��~ �~P�L$Dv(��	f/�v(�f/�v(��	f/�v(�f/�wf/�v(��(ġ|A�$�T$�\$�@�$�@HQ�t$<�L$<�Ѓ�0���̡|A�@H��0  ���������������������������������̡|A�@H���  ��|A�@H���  ���t$,�|A�t$,�@H�t$,���  �t$,�t$,�t$,�t$,�t$,�t$,�t$,�t$,Q�Ѓ�0�, ��������������t$,�|A�t$,�@H�t$,���  �t$,�t$,�t$,�t$,�t$,�t$,�t$,�t$,Q�Ѓ�0�, ������������̡|AQ�@H��,  �Ѓ������������̡|A�t$�@HQ��X  �Ѓ�� ����̡|AQ�@H��\  �Ѓ������������̡|AQ�@H�t$���   �t$�Ѓ�� �SUV�t$W�|$3ҋ���ƃ�t��    ��B��u��PSWU�L$$��  �� ~%��   VWU�L$ �q  SVU�L$ �  _^][� ;�tSWU�L$ �N  _^][� �������V���v���|A�@l�@�Ѓ��D$t	V�������^� �������������̃�U�l$����   �L$��S�V+���F�Y�W�6�<��t$�D$(�|$�\$��\$�|$�D$(�d$ ��~N�����t$�\$�D$(�&�G���S����GM�C�|$��W��~g�L$$����9l$(���    ���G���;�}�;H}G���;�t$�L$$�u������s��H�K�?;͋L$$��p~��t$�M���_^[]��� ��̋T$U�l$��+����� ~PU�t$�����]� SVW�]��    ��;�t(�;H�}�p�ыH���H��H�P��p����;�u܋T$��;�u�_^[]� ����QS�\$W�|$��+ǃ���L$=   ��   U�l$ V��tv�7��+����+����K��Ǎ�M�T$ ;�}9T$ |��;��;�}���9T$ L��L$PSW�t$$�   �L$US��V�t$$�v�����+������   �^]_[Y� �L$SW�t$ �����^]_[Y� ��������S�\$V�t$;�t4UW��F���;}�n����
�H�@��J�R�;8|�:�j��;�u�_]^[� ��������̋D$S�\$VW�|$�����9|���I ��;|�;�s$���p��O�H��w;�u����;�uǋ���_^[� �����������U�������  V��MW�t$D��u'�E�~f� �~Ff�@�~Ff�@_^��]� �}���^�G0�V�o �Y�f(��Y�f(��Y��X'�FP�Xw�X��GH�Y��X��d$�d$ �g8(��Y��X��GP�Y��X��t$�t$(�w((��Y��D$8���G@�XO�Y��X��GX�Y��X��L$8�L$0����  �$�<(�f �V�^((��YG0(��Y��Y�E�X�(��YGH�Y�j �X��G8�Y�j ����$   �X��GP�Y��X��G@�Y���$(  �X��GX�Y��X��D$ ��$h  �D$0��$p  �D$P��$x  �@�D$� �$��$   P��$l  P��$  P��$<  躮  ��  �f �V�^((��YG0(��YύD$8P�E�X�(��YGH���X�(��Y��Y���$�   (��YO8�Yg@�X�(��YGP�Y_X�X��X��D$��$�  �D$,��$�  �D$L��$�  �@�D$� �$��$�   P�X㍄$�  P��$�  P��$�   ��$�   �>�  �|$8 �~ f�D$ �~@f�D$(�~@f�D$0��
  �O�Y�f�G0�^�X�Y��w8�(�M�X��GH�YÍ�$�   P��$D  �X�(��Y��gX��$�   �O �YP�XO�X��GP�Y��_@�X�(��YF��$�   (��Y�XO�X�(��YF�X���XF��$�   �N�XN �D$�Y|$�L$ �N�XN(�X�Yt$ �Y\$ �L$�O�Y��G0�YD$ �X�Yd$�X��X��GH�YD$�X��X��GP�YD$��$�  ��$p  �O �YL$�XO�X��X���$x  �  ����$h  P��$4  �MP�  � �\�D$`�@�\F�D$h�@�\F�D$`P��$t  P�D$x�  �`�H�(�t$L�wW��Y�f(��Y��\�f(��\��Y��V�L$P��\��Y��\$X�^�g(�X7f(��YG0�l$`(��Yo �X��GH�Y��Xo�M�Y��X�(��YG8�Xg����$�  �X��GP�Y�P��$  P�X��G@�Y��t$�l$��$�  �X��GX�Y���$�  �X��d$ ��$�  �H  �P�H�XT$P�XL$X�D$H�X �M��$8  P��$�  P��$@  ��$H  ��$P  �U  � �\D$�D$`�@�\D$�D$h�@�\D$�D$`P��$d  P�D$x��  �~ ��O�f�^f�D$P�~@f�D$X�~@�Y�f�D$`(��YG0�X�E�M���X��GH�Y�j j ���X�(��YG8��$�   (��YO �XO�X��GP�Y��X��G@�Y���$�   �O(�Y��XO�X��GX�Y��X��@�D$� �$�D$`P��$�   P��$0  P��$�   �&�  �7  �U�Bf. ���D{R��$,  �  ��D$ P�D$�B��$\  P�D$�  �@�L$��$�   ��$�   �L$P��$�   ��$�   ��$�  �  �f �V�G0�^(�Y�(��YʋEj ���X��GH�Y��X��G8�Y���$  (��Y��X��GP�Y��X��G@�Y��gX��$  (��Y��V8�X�(��Y��_0�Y��X��F0�Y��Y���$  �X?�N@�Xo�Y��G@�X��_H�Xw�Y��Y��Y��X��_8�Y��X��@�D$� �X��_P�Y��$��$  P�X��X�$8  P��$�  P��$@  ��$H  ��$P  豧  �~�\$ �\^0�~H�L$(�~P�\$�\N8�\V@f(��Y��L$(��Y��T$�X�(��Y��X��o�  f(�W�f.ʟ��Dz
f(�f(��*���^��T$�L$�\$�Y��Y��Y��FH�Y��Y��Y��XV0�XN8�X^@f�T$ f�L$(f�\$0�  �F0�V8�_0�N@�Y��Y��Y��X?�Y��G@�Xw�X��_H�Xo�Y��Y��Y��X��_P�X��GX�X��Y��Y�j�X�D$|�X�P��$�   ��$�   ��$�   讥  �\$�D$�YFHf. �D$���Dz��L$�V0�O�f8�^@�Y�(��YG0�X�M��$�  P��$�  �X�(��YGHP�X�(��YG8��$�  (��YO �XO�X�(��YGP�X��G@�Y���$�  �O(�Y��XO�X��GX�Y��X���$�  �y  �M��\�I�\H�T$f(��Y��L$(��Y�W��X�(��Y��X��.�  �d$f(�f/�vf(��f(�W�f.џ��Dz
f(�f(��'���^��T$�\$�Y��Y��Y�(��Y��Y��Y��^��f�T$(f�\$0f�L$8�,$��  ���\$�D$菮  �YD$�V0�O�f8fW0�^@�Y��D$0f(��YG0�X�M��$�  P��$  �X�f(��YGHP�X�f(��YG8��$�  (��YO �XO�X�f(��YGP�X��G@�Y���$�  �O(�Y��XO�X��GX�Y��X���$�  ��  �P�H� �XT$(�XL$0�XD$ ��$�  P��$�  ��$�  ��$�  ��$L  �MP��  �~ f�D$ �~@f�D$(�~@f�D$0��$x  WP�L
  �d$(�\$0�T$8�ȋE�I�A0�Y��YÃ��X	_^�X��AH�Y��X��A8�Y���I �Y��XI�X��AP�Y��X��A@�Y��H�I(�Y��XI�X��AX�Y��X��H��]� ���/!�!�#� �������������U������   �}SVW�L$t�   _^[��]� �}�W�Px�D$��t�|A�]�@HS��   W�Ћ|A�u�Id�D$�I<�ы��D$|j/P�1  ��$�   jP�1  �|AV�@dW�@pS�Ѓ�(3��|Aj �@d��$�   �@��t�L$tQS��3���9t$��   �L$3�;���;���   �L$W���T$RV�uf�D$$f�D$,f�D$4f�D$<f�D$Df�D$Lf�D$Tf�D$\f�D$d���D$l�D$t    �P|�|$h�t�|Aj �@dj���   �L$ QS�Ѓ��L$F;t$�]���G��� ���_^�   [��]� �������������̸   � ��������U�������   �ESVW��t���_^[��]� �|A�L$�@HQ�M�@,�Ћ���   ��$�   �}W���D$����3��Px���z  �W��L$Qf�D$f�D$f�D$$f�D$,f�D$4f�D$<f�D$Df�D$Lf�D$T��VW���D$d�D$l    �P|�|$`��  �d$��$�   �\$��$�   �T$ �Y��Y��u�X�$�   �|A�u�L$xQ�X���$�   �Y��u�X���$�   �Y���$�   ��$�   �Y��X�$�   �X���$�   �Y��X���$�   �Y���$�   ��$�   �Y��X�$�   �X���$�   �Y��X���$�   �@d�@�Ѓ���t
�E�t$t�W��F�Rx;�������D$_^[��]� ����U������4  �|AS�@HV�@$�L$�MW�Ћ|A�M�RH�؋R<��$�   P���#�S�[f(̹   ���|$��YL$(�|$8f(��YD$@�XL$�t$P�l$h�X�f(��YD$X�X�f(��YD$H�Y���$�   f(��YL$0�Y��XL$�Xd$ �X�f(��YD$`�X��S(�Y��X��X��[ ��$�   f(��YD$@��$�   �cf(��YL$(�X�f(��YD$X�X�f(��YD$H�Y���$�   f(��YL$0�Y��X�f(��YD$`�X��Y��X��X���$�   ��$�   �[8�c0�S@f(��YL$(f(��YD$@�|A�uj �X�f(��YD$\V�X�f(��YD$P�Y���$   f(��YL$8�Y��X�f(��YD$h�X��[P�Y��X�f(��YD$H�X��SX��$  ��$  �cHf(��YL$0Ǆ$�       �X�f(��YD$`�X�f(��YD$P�Y���$  f(��YL$8�Y��X�f(��YD$h�X��Y��X�W�f�D$xfք$�   fք$�   fք$�   fք$�   fք$�   fք$�   fք$�   fք$�   ���X���$�   �@@��$   �@8��$(  �Ћ}����L$pQWV���R|�u�\$��$�   �3P�u��$4  P��$�   �N����~ �L$pQ����W�uf��~@f�A�~@f�A�����   _^�   [��]� ��������������3�� �����������3�� ������������ �������������3�� ����������̸   �$ ��������� �������������3�� ������������ �������������3�� ������������ ��������������$ ������������̡|A�L$�@��   �@<�Ѕ�t#j ��$8  ��$,  �P�������u��   �Sh   �D$j P�8�  ��$<  j ��$L  �D$��$T  S��$P  P�   ��$�   ����5E���$�   ��$�   �� ��5E���$�   ��$�   �À��5E���$�   ��$�   ��5��E�h   ��$�   �D$,P��$X  Ǆ$�   �5��$X  j��#  ��8[��   ���������������V�t$W�t$ �|$�t$V�t$�t$$W�_1�������   Ǉ�   �5Ǉ�   �5Ǉ�   �5Ǉ�   �5Ǉ�   �5Ǉ�   �5Ǉ�   �5Ǉ�   �5_^����U�������   VW�M�qX�I8�y(�A@�YAP�Y�f(��YQP�D$X�L$H�\��A �D$`�Y�f(��T$8�Q �YQ@�\��D$h(��YA8�T$ �L$0�D$(��Q0�\��A�Y��Y�W��|$(�\$@�X��AH�Y��d$P�X���f.џ��DzD�Ef�f�@f�H0f�HHf�Hf�H f�@8f�HPf�Hf�H(f�H@f�@X_^��]��^��y�D$�A(��Y�(��Yq@(��Ya8�(��YYP(��Yy �\��d$(��\��d$h�YA0�\d$8�YIH�\t$�\��i�X��D$X�\D$H�Y��Y��Y��Y��X��YL$�L$p�I�YL$((��\��\��YAH�Yy0�X��X��\$�Y��D$x�D$�\D$ �Y��QH(��YI@�X��D$0�Y��X��y0��$�   �D$@�Y��Y���$�   �D$P�Y���$�   ��$�   (��YAX�\�(��YA(�Y���$�   (��YIX�\��Y���$�   (��YI((��YA@�E�t$p���\�(��YA8�YT$`�Y���$�   (��YIP�Y|$`�\�(��Yi8�YAP�Y��\��\й   ��$�   �Y��Y���$�   ��$�   �_^��]����U����QV�u�V��^(��Y��Y��X�(��Y��X�脟  f(�W�f.џ��D�Ez��H�H^��]����^���Y���N�Y��H�N�Y�^�H��]Ë�`D��`H��`L��`P��`T��`X��`\��``��`d��`h��`l��`p��`t��������L$f/�r���f/�r� �(�蜞  �D$�D$�̡|A���@h�t$ �@0Q�L$Q�ЋL$(�~ f��~@f�A�~@f�A����$� �������������̡|A���@h�t$ �@8Q�L$Q�ЋL$(�~ f��~@f�A�~@f�A����$� �������������̡|A���@h�t$ �@,Q�L$Q�ЋL$(�~ f��~@f�A�~@f�A����$� �������������̋D$V�0W�9;�t_3�^� �P��u��u9pu9qu��u�9yu�_�B^� S�Y��u!��u9yu��u2��u.9pu)[_�   ^� ��t��t;�u�P��t�A��t�;�t�[_3�^� �������t$�g������@� ���������������VhhAj\hD ��茗  ����t�@\��tV�Ѓ���^�����VhhAj\hD ���\�  ����t3�@\��t,V��hhAjxhD �:�  ����t�@x��t
V�t$�Ѓ���^� �����������̃�VhhAj\hD �����  ����tL�@\��tEV�ЋD$hhAjdhD �D$�D$    �D$    迖  ����t�@d��t�L$QV�Ѓ���^��� �������������VhhAj\hD ���|�  ����t3�@\��t,V��hhAjdhD �Z�  ����t�@d��t
�t$V�Ѓ���^� ������������VhhAj\hD ����  ����t\�@\��tUV��hhAjdhD ���  ����t�@d��t
�t$V�Ѓ�hhAjhhD �ѕ  ����t�@h��t
�t$V�Ѓ���^� ���VhhAj\hD ��蜕  ������   �@\��t~V��hhAjdhD �v�  ����t�@d��t
�t$V�Ѓ�hhAjhhD �M�  ����t�@h��t
�t$V�Ѓ�hhAjhhD �$�  ����t�@h��t
�t$V�Ѓ���^� ������VhhAj`hD ����  ����t�@`��tV�Ѓ�^�������VhhAjdhD ��輔  ����t�@d��t
�t$V�Ѓ�^� VhhAjhhD ��茔  ����t�@h��t
�t$V�Ѓ�^� VhhAjlhD ���\�  ����t�@l��tV�Ѓ�^�������VhhAjphD ���,�  ����t�@p��t�t$V�Ѓ�^� �lA^� �������VhhAjxhD ����  ����t�@x��t
V�t$�Ѓ���^� ��������������VhhAj|hD ��謓  ����t�@|��tV�t$�Ѓ�^� 3�^� ����������VhhAj|hD ���l�  ����t�@|��tV�t$�Ѓ����@^� �   ^� ��j�h��d�    P��V�8A3�P�D$d�    ��hhAjthD �D$    ��  ����tu�@t��tn�t$(�L$VQ�Ѓ��t$$P���D$    �`���hhAj`hD �D$   �D$( 貒  ����tv�H`��to�D$P�у��ƋL$d�    Y^��� hhAj\hD �t�  �t$0����t4�@\��t-V��hhAjdhD �N�  ����t�@d��thlAV�Ѓ��ƋL$d�    Y^��� VhhAh�   hD ���	�  ����t���   ��t�t$V�Ѓ�^� 3�^� ����VhhAh�   hD ���ɑ  ����t���   ��t�t$V�Ѓ�^� 3�^� ����VW��3����$    �hhAjphD ��  ����t�@p��t	VW�Ѓ���lA�8 tF��_��^�������SU�l$V��3�W�d$ hhAjphD �/�  ����t�@p��t	VS�Ѓ���lA�8 tnhhAjphD ���  ����t�@p��tVU�Ѓ�����lAhhAjphD �ΐ  ����t�@p��t	VS�Ѓ���lAW���Z�����tF�`����D$_��t�0��~=hhAjphD 耐  ����t�@p��t	VS�Ѓ���lA�8 u^]�   [� ^]3�[� �����������̃�VhhAh�   hD ���&�  ����t?���   ��t5�t$�L$VQ��hhAj`hD ���  ����t�@`��t
�L$Q�Ѓ���^��� �������j�h�d�    P��V�8A3�P�D$d�    hhAh�   hD �D$    萏  ����ty���   ��to�t$,�L$�t$,Q�Ѓ��t$$P���D$    �����hhAj`hD �D$   �D$( �;�  ����ts�H`��tl�D$P�у��ƋL$d�    Y^���hhAj\hD ���  �t$0����t3�@\��t,V��hhAjxhD �َ  ����t�@x��t
V�t$,�Ѓ��ƋL$d�    Y^����������������̋���������������hhAjhD ��  ����t	�@��t��3��������������V�t$�> t+hhAjhD �E�  ����t�@��tV�Ѓ��    ^���������̃|$ W��t1hhAjhD ��  ����t�@��t�t$�t$W�Ѓ�_� 3�_� ���������������VhhAjhD ��輍  ����t�@��t�t$V�Ѓ�^� 3�^� ����������VhhAjhD ���|�  ����t�@��t�t$V�Ѓ�^� 3�^� ����������VhhAj hD ���<�  ����t�@ ��tV�Ѓ�^�3�^���VhhAj$hD ����  ����t�@$��tV�Ѓ�^�3�^���VhhAj(hD ���܌  ����t�@(��t�t$�t$�t$V�Ѓ�^� 3�^� ��VhhAj,hD ��蜌  ����t�@,��t�t$�t$V�Ѓ�^� 3�^� ������VhhAj(hD ���\�  ����t�@0��t�t$�t$�t$V�Ѓ�^� 3�^� ��VhhAj4hD ����  ����t�@4��tV�Ѓ�^�3�^���VhhAj8hD ����  ����t!�@8��t�t$�t$�t$�t$V�Ѓ�^� 3�^� ��������������VhhAj<hD ��蜋  ����t�@<��t
�t$V�Ѓ�^� VhhAh�   hD ���i�  ����u^� �t$���   V�Ѓ�^� ����������VhhAh�   hD ���)�  ����u^� �t$���   V�Ѓ�^� ����������VhhAh�   hD ����  ����u^� �t$���   V�Ѓ�^� ����������VhhAh�   hD ��詊  ����t�t$���   �t$�t$V�Ѓ�^� ������VhhAjDhD ���l�  ����t�@D��tV�Ѓ�^�3�^���VhhAjHhD ���<�  ����t�t$�@HV�Ѓ�^� ����VhhAjLhD ����  ����u^� �t$�@LV�Ѓ�^� VhhAjPhD ���܉  ����u^� �t$�@P�t$V�Ѓ�^� ������������VhhAh�   hD ��虉  ����u^� �t$���   �t$�t$V�Ѓ�^� ��VhhAh�   hD ���Y�  ����u^� �t$���   �t$�t$�t$�t$V�Ѓ�^� ����������VhhAjThD ����  ����u^Ë@TV�Ѓ�^���������VhhAjXhD ���܈  ����t�t$�@XV�Ѓ�^� ����j�hI�d�    P��V�8A3�P�D$ d�    ��hhAh�   hD �D$    �~�  ����t~���   ��tt�t$4�L$Q���Ћt$0P���D$,   �����hhAj`hD �D$   �D$4 �.�  ������   �H`����   �D$P�у��ƋL$ d�    Y^��$� hhAj\hD �D$     �D$$    �D$(    �Ї  �t$<����t4�@\��t-V��hhAjdhD 誇  ����t�@d��t�L$QV�Ѓ��ƋL$ d�    Y^��$� ������������VhhAh�   hD ���Y�  ����t���   ��t�t$���t$�t$��^� 3�^� ��������������VhhAh�   hD ���	�  ����t���   ��t�t$����^� 3�^� ������VhhAh�   hD ���Ɇ  ����t���   ��t�t$����^� 3�^� ������VhhAh�   hD ��艆  ����t���   ��t�t$����^� 3�^� ������VhhAh�   hD ���I�  ����t���   ��t��^��3�^����������������VhhAh�   hD ���	�  ����t���   ��t�t$���t$�t$��^� 3�^� ��������������VhhAh�   hD ��蹅  ����t���   ��t�t$����^� ������������VhhAh�   hD ���y�  ����t���   ��t�t$���t$�t$��^� 3�^� ��������������VhhAh�   hD ���)�  ����t���   ��t��^��3�^����������������hhAjhD ��  ����t	�@��t��3��������������j�h��d�    P��VW�8A3�P�D$ d�    hhAh�   hD �D$    菄  ����u)�|A�t$0�HV�I�у��ƋL$ d�    Y_^�� ��t$4���   �L$Q�Ћ��|A�|$8�IW�I�D$4   �ѡ|AW�@V�@�Ћ|A�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� ������������hhA�t$hD �̓  ������������hxAjh�f 诃  ����t	�@��t�����������������j�h��d�    PQV�8A3�P�D$d�    hxAjh�f �D$     �U�  ������t9�~ t3�t$L�D$$�t$L�t$L�t$L�t$L����P�����t$L�F�Ѓ�4�������L$ �D$�����o����ƋL$d�    Y^���������������hxAjh�f �ς  ����t	�@��t��3��������������hxAjh�f 蟂  ����t	�@��t��3��������������hxA�t$h�f �m�  �����������̋D$�|A� ����̡|AQ���   �@X�Ћȃ���u� �|A�t$�@|�t$�@Q�Ѓ�� ������̡|AQ���   �@X�Ћȃ���u� �|A�t$�@|�t$�@8Q�Ѓ�� ������̋T$V��j ��|Aj �@j �@R�Ѓ��F��^� ������̡|AV�@j �@j ��j �6�Ѓ��F^�V��N��u3�^� �|AQ�t$�@�t$�@�6�Ѓ��F�   ^� ��������̋D$HV����   �$�,O�   ^á�A@��A��uU�t$������=�6  }�����^Ët$��t�jh@jmj���������t	���S����3���A��tV�������   ^��t$�t$�J����������H^�^������Au.�����%����5�A��t�������V��������A    �   ^Ã��^Ð]N�N�NVN&O�N�������������L$u�D$��A�D$��A�   � �|AV�@j �@j����Ћ�^��������̡|AV�@j �t$�@���Ћ�^� ���̡|AV�@�t$�@j����Ћ�^� ���̡|A�@�@����̡|AV�@j ���   ��L$j V�Ћ�^� �������������̡|A�t$�@Q�@�Ѓ�� �������̡|A�t$�@Q�@�Ѓ����@� ��̡|Ah#  �t$�@�t$�@l��� ��̡|AhF  �t$�@�t$�@l��� ��̡|A�t$�@�@t�Ћ|AP���   �@X�Ѓ�� ������̡|A�t$�@�@t�Ћ|A�t$�Ћ��   R�@`�Ѓ�� ̡|A�t$�@���   �Ћȅ�u� �|AQ���   �@�Ѓ�� �����������̡|A�@���   ��|A���   �AP���   ��Y�������̡|A�t$�@8Q�@D�Ѓ�� �������̡|A�@8�@<����̡|AV�@8�t$�@@�6�Ѓ��    ^���t$�|A�t$�@8�t$�@�t$�t$�t$Q�Ѓ�� �����t$�|A�t$�@8�t$�@�t$�t$Q�Ѓ�� �������̡|A�@8� �����̡|AV�@8�t$�@�6�Ѓ��    ^���t$�|A�t$�@8�t$�@Q�Ѓ�� �|A�t$�@8�t$�@Q�Ѓ�� ���̡|AQ�@8�@�Ѓ���������������̡|A�t$�@8Q�@ �Ѓ�� ���������t$�|A�t$�@8�t$�@$�t$�t$Q�Ѓ�� �������̡|A�t$�@8�t$�@(Q�Ѓ�� �����t$�|A�t$�@8�t$�@,Q�Ѓ�� �t$�|A�t$�@8�t$�@Q�Ѓ�� �|A�t$�@8�t$�@0Q�Ѓ�� �����t$�|A�t$�@8�t$�@4Q�Ѓ�� �|A�t$�@8Q�@8�Ѓ�� �������̋L$�|A�P�APP�A@P�A0P�A P�AP���   Q�t$�Ѓ����������������̡|A�@���   ��|A�@���  ��|A�@�@,����̡|A�@���  ��j�h��d�    PQV�8A3�P�D$d�    �D$    �|A�t$�@V�@�D$    �Ћ|AV�I�D$    �I8�D$   �у��ƋL$d�    Y^���������̡|A�@�@<����̡|A�@�@@����̡|A�@�@D����̡|A�@�@H����̡|A�@�@L����̡|A�@�@P����̡|A�@��<  ��|A�@��,  ���t$�|A�t$�@�t$���   �t$�t$h�6  �Ѓ����̡|A�@�@�����j�h�d�    P�� �8A3�P�D$$d�    �|A�L$�@Q�@�С|Aj �@j��@�L$h�Q���t$H�D$P�D$0P�D$L    �5����|A�L$$�@Q�@�D$P�С|A�L$8�@Q�@�С|A�L$<�@Q�@�D$X�����Ѓ�,�L$$d�    Y��,���������������̡|A�@���  ��|A�@��8  ��j�hL�d�    P��VW�8A3�P�D$ d�    �D$    �|A�L$�@Q��  �Ћ��|A�|$4�IW�I�D$0   �ѡ|AW�@V�@�Ћ|A�D$ �IP�I�D$    �D$< �у��ǋL$ d�    Y_^�� ������������j�h��d�    P��VW�8A3�P�D$ d�    �D$    �|A�L$�@Q��  �Ћ��|A�|$4�IW�I�D$0   �ѡ|AW�@V�@�Ћ|A�D$ �IP�I�D$    �D$< �у��ǋL$ d�    Y_^�� �����������̡|A�@��x  ��|A�@��|  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@�@T����̡|A�@�@X����̡|A�@�@\����̡|A�@�@`����̡|A�@���  ��|A�@�@d����̡|A�@�@h����̡|A�@�@l����̡|A�@�@p����̡|A�@�@t����̡|A�@��D  ��|A�@��  ��|A�@�@x����̡|A�@��@  ��j�h��d�    PQV�8A3�P�D$d�    �D$    �t$���D$    ������|AV�I�t$$�I|�D$    �D$   �у��ƋL$d�    Y^������������̡|A�@���   ��|A�@��d  ��|A�@��h  ��|A�@���  ��|A�@���   ��j�h��d�    PQV�8A3�P�D$d�    �D$    �t$���D$    �s����|AV�I�D$    ���   �D$   �у��ƋL$d�    Y^�������������̡|A�@��`  ��|A�@��  ��|A���@�t$ ���   �L$Q�ЋL$$�~ f��~@f�A�~@f�A���� ��������������̡|A�@���  ���t$�D$�|A���@�D$�D$���   �$�t$�Ѓ�����������̡|A�@���   ��|A�@���   ��|A�@���  ��|A�@���  ��|A�@��   ��|A�@��  ��|A�@��l  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@���  ��j�h$�d�    P��VW�8A3�P�D$ d�    �t$4�D$    �|A�L$�@Q���  �Ћ��|A�|$8�IW�I�D$4   �ѡ|AW�@V�@�Ћ|A�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� ��������j�h`�d�    P��VW�8A3�P�D$ d�    �t$4�D$    �|A�L$�@Q���  �Ћ��|A�|$8�IW�I�D$4   �ѡ|AW�@V�@�Ћ|A�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� �������̡|A�@���  ��|A�@���  �����|A�T$�@R���   �T$R�T$RQ�����#D$���̃��|A�T$�@R���   �T$R�T$RQ�����#D$���̃��|A�$�@R���   �T$R�T$RQ�����#D$����̡|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@��  ��|A�@��\  ��j�h��d�    P�� �8A3�P�D$$d�    �t$8�D$    �|A�L$�@Q��t  �Ѓ��t$4���D$0   ������L$�D$   �D$, � ����D$4�L$$d�    Y��,������������̡|A�@��H  ��|A�@��T  ��|A�@��p  ��|A�@��8  ����  �8A3ĉ�$   ��$  P��$  �D$h   P�\ ����x	=�  |'��|Ah��@hH  ��0  �Ѓ�Ƅ$�   �|A�$�@Q��4  h��Ћ�$  ��3��p  ��  �������������������������t$$�D$�t$$�P�t$$�|A�t$$�@0�t$$���   �t$$�t$$�t$$RQ�Ѓ�(�$ ��t$$�D$�t$$�P�t$$�|A�t$$�@0�t$$���   �t$$�t$$�t$$RQ�Ѓ�(�$ ��t$$�|A�t$$�@0�t$$���   �t$$�t$$�t$$�t$$�t$$�t$$Q�Ѓ�(�$ ����̡|AQ�@0���   �Ѓ������������̡|A�t$�@0�t$���   Q�Ѓ�� ��t$�|A�t$�@0�t$���   �t$Q�Ѓ�� ��������̡|AQ�@0���   �Ѓ��������������t$�|A�t$�@0�t$���   �t$Q�Ѓ�� ��������̡|A�@0���   ��|AV�@0�t$���   �6�Ѓ��    ^���������������j�h��d�    P��V�8A3�P�D$d�    �t$8�D$    �|A�t$8�@�t$8��X  �L$Q�ЋЋt$<j �    �F    �|AR���   V�@�D$@   �Ћ|A�D$(���   P�	�D$(   �D$D �у� �ƋL$d�    Y^�� ������������j�h�d�    P��(V�8A3�P�D$0d�    hLGOg�L$ �D$    �����j P�D$hicMCP�D$H   ��������L$�D$8�����|A�L$���   Q�@T�Ѓ���u�L$@�����"�|A�L$���   Q�@T�ЋL$D��P�����|A�D$���   P�	�D$   �D$< �ыD$D���L$0d�    Y^��4��������̡|A�@���  ��|A�@���  ��|A�@���  ��j�hT�d�    P��VW�8A3�P�D$ d�    j �t$D�D$    �t$D�|A�t$D�@�t$D��t  �L$$Q�Ћ��|A�|$H�IW�I�D$D   �ѡ|AW�@V�@�Ћ|A�D$4�IP�I�D$4   �D$P �у�(�ǋL$ d�    Y_^�� ����������j�h��d�    P��V�8A3�P�D$d�    �t$<�D$    �t$<�|A�t$<�@�t$<���  �L$Q�ЋЋt$@j �    �F    �|AR���   V�@�D$D   �Ћ|A�D$,���   P�	�D$,   �D$H �у�$�ƋL$d�    Y^�� ��������j�h��d�    P��$�8A3�P�D$(d�    �|A�@��p  �Ѕ���   h���L$�G����|A�t$8�@h���@4�L$�D$8    �С|A�t$<�@h���@4�L$��j �D$P�D$hicMCP�����|A�L$���   Q� �Ѓ��L$�D$0���������L$(d�    Y��0��������������j�h��d�    P��(VW�8A3�P�D$4d�    �D$    �|A�@��p  �Ѕ�u)�|A�t$D�HV�I�у��ƋL$4d�    Y_^��4�h!���L$$�8����|A�t$H�@h!���@4�L$(�D$D   ��j �D$$P�D$hicMCP����P�|A�D$P���   �@H�Ћ|A�|$X�IW�I���ы|AW�AV�@�Ћ|A�D$0���   P�	�D$0   �D$`�у�$�L$ �D$< ������ǋL$4d�    Y_^��4��������������j�h;�d�    P��(VW�8A3�P�D$4d�    �D$    �|A�@��p  �Ѕ�u)�|A�t$D�HV�I�у��ƋL$4d�    Y_^��4�h����L$$������|A�t$H�@h����@4�L$(�D$D   ��j �D$$P�D$hicMCP�����P�|A�D$P���   �@H�Ћ|A�|$X�IW�I���ы|AW�AV�@�Ћ|A�D$0���   P�	�D$0   �D$`�у�$�L$ �D$< �����ǋL$4d�    Y_^��4��������������j�hf�d�    P��$V�8A3�P�D$,d�    �|A�@��p  �Ѕ�u�L$,d�    Y^��0�h#���L$������|A�t$<�@h#���@4�L$ �D$<    ��j �D$P�D$hicMCP����P�|A�D$H���   �@8�Ћ|A�����   �D$�	P�D$L �у��L$�D$4���������ƋL$,d�    Y^��0��������j�h��d�    P��$V�8A3�P�D$,d�    �|A�@��p  �Ѕ�u�L$,d�    Y^��0�hs���L$������|A�t$<�@hs���@4�L$ �D$<    ��j �D$P�D$hicMCP�����P�|A�D$H���   �@8�Ћ|A�����   �D$�	P�D$L �у��L$�D$4���������ƋL$,d�    Y^��0�������̡|A�@���  ��|A�@���  ��|A�@��@  ��V�t$���t�|AQ�@��D  �Ѓ��    ^���������̡|A�@��H  ��|A�@��L  ��|A�@��P  ��|A�@��T  ��|A�@��X  ��|A�@��\  ��|A�@��d  ��|A�@��h  ��|A�@��l  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@��P  ��|A�@���  ��j�h��d�    P���8A3�P�D$d�    �t$0�D$    �|A�L$�@Q���  �Ѓ��L$,P�D$(   ������L$�D$   �D$$ ������D$,�L$d�    Y��$�������������̡|A�@���  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@���  ��|A�@��l  ��|A�@���  ��|A�@���  ��|A�@��$  ��|A�@��(  ��|A�@��,  ��|A�@��0  ��|A�@��<  ��|A�@��  ��|A�@��`  ��|A�@��\  ���� ��V���.�vf(�fT�	f/�f(�fT�	�T$�L$�L$�-  f/��#  �X	f/�vFf/�v@�,��,���   ��$    ������ʅ�u�fn�����^��^��.�v^�� �f/�v(��(��h	�^��%�f/�v4(��Y��Y��Y��D$(��Y��.�v(��L$�L$f/�v(��D$�D$�f��D$�D$�f  �\$�D$f/P	�L$�L$�D$�D$s���^���F�^��F^�� �W�����F^�� �����������������D$�`	f/�V��w�p	f/�v(��Y����XP	�D$�D$�$�e  ��������F�������^� ���̃��L$�T$3�W�f/�fT�	�XP	��3�f/�V����3��L$�D$;������$�L$�=e  ��D$ fT�	�D$ �XP	�D$ �D$ �$�e  ���\$ �D$ ��f/��Fv'�|Ah��@j��0  �������F�|$ u�fW0���������^��� ������������D$��f/�V���Fv'�|Ah��@j,��0  �������F^� ���������U�����M����<f/�V��v'�|Ah$	�@j5��0  �������M��Y����D$8�D$8�$��c  �\$8�F�$��c  �D$8�\$@�^D$@�D$@�D$@�$�c  ��E�$�c  ���^�������^��]� ����������̋L$��`������̋L$��`�������V��hpt��	�F    �|AV�@PhPq� h@q�Ѓ��F��^����������̃y ��	u�|A�q�@P�@��Y��̋I��u3�� �|Aj �t$�@P�t$�@Q�Ѓ�� �����̋I��t�|A�t$�@PQ�@�Ѓ�� ̋I��t�|A�t$�@PQ�@�Ѓ�� ��    �A    ���V����t&�|AQ�@P�@L�С|A�6�@P�@<�Ѓ��    ^����������������SUVW�����t�|AQ�@P�@<�Ѓ��    �G    �\$�l$hptS�o�|AhPq�@Ph@q�@8U�t$(�Ѓ�3����~D���x u�@   �|A�HP���p�A�Ѓ��|AV�@P�7�@@�Ћ�F���A;�|�3�9_^]��[� �������������t$�D$�t$�p�,���� ���������SVW��3�9w~>�\$�|AV�@P�7�@@�ЋЃ���t,�|Aj �APS�@jR�Ѓ���tF;w|�_^�   [� �|A�7�@P�@L�Ѓ�3�_^[� ̡|A�1�@P�@D�Ѓ��������������̡|A�1�@P�@H��Y���������������̡|A�1�@P�@L��Y���������������̡|A�@P�@P����̡|A�@P�@T����̡|A�@P���   ��|A�@P���   ���L$��`�������V��~ ��	u�|A�v�@P�@�Ѓ��D$t	V聩������^� ��������3��������������̡|AQ�@L���   �Ѓ������������̡|A�t$�@L�t$���   Q�Ѓ�� ̡|AV�@L�񋀠   V�Ћȡ|A����u�@LQ�t$���   V�Ѓ�^� ���   �@P�Ћ|AP���   �L$�BH��^� ̡|AQ�@L��(  �Ѓ������������̡|A�t$�@L�t$��,  Q�Ѓ�� ̡|A�@L� �����̡|AV�@@�t$�@�6�Ѓ��    ^�̡|A�@L���   ��|AV�@@�t$�@�6�Ѓ��    ^��j�h�d�    P���8A3�P�D$d�    �t$0�D$    �|AQ�@L�L$�@Q�Ѓ��L$,P�D$(   �I����L$�D$   �D$$ �S����D$,�L$d�    Y��$� ������������̡|A�t$�@L�t$�@Q�Ѓ�� ���̡|A�t$�@LQ���   �Ѓ�� ����̡|AQ�@L�@�Ѓ���������������̡|AQ�@L�@�Ѓ���������������̡|AQ�@L�@�Ѓ�����������������t$�|A�t$�@L�t$�@ Q�Ѓ�� �|A�t$�@LQ��4  �Ѓ�� ������t$�|A�t$�@L�t$�@$Q�Ѓ�� �t$�|A�t$�@L�t$�@(�t$Q�Ѓ�� �����������̡|AQ�@L�@,�Ѓ���������������̡|AQ�@L�@0�Ѓ���������������̡|AQ�@L�@4�Ѓ���������������̡|Aj �@LQ�@8�Ѓ�������������̡|A�t$�@L�t$��  Q�Ѓ�� ̡|A�@L���   ��|A�@L���   ��|A�@L��l  ��|A�@L���   ��|A�@L���   ��|A�@L���   ��|A�@L���   ��|A�@L���   ��|A�@L���   ��|A�t$�@LQ�@<�Ѓ�� �������̡|A�@L���   ��|AQ�@L�@��Yá|A�t$�@L�t$�@@Q�Ѓ�� ���̡|Aj �@L�t$�@DQ�Ѓ�� �����̡|Aj�@L�t$�@DQ�Ѓ�� �����̡|Aj �@L�t$�@HQ�Ѓ�� �����̡|Aj�@L�t$�@HQ�Ѓ�� �����̡|AQ�@L���   �Ѓ�������������j�hE�d�    P���8A3�P�D$d�    �t$0�D$    �|AQ�@L�L$��  Q�Ѓ��L$,P�D$(   �V����L$�D$   �D$$ �`����D$,�L$d�    Y��$� ����������j�hp�d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �����j �D$$P�D$P���D$D��������L$���D$8 �`�����t3���|A�L$ ���   Q�@8�Ѓ����|A�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h��d�    P��$V�8A3�P�D$,d�    ���D$   �D$$   �D$P�L$�D$8    �D$�  �D$    �D$    ����j�D$ P�D$P���D$@�����L$�D$4 �v����|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0�������j�h��d�    P��(SV�8A3�P�D$4d�    ���D$    �D$$    �D$,    �D$P�L$�D$@   �D$�  �D$     �D$$    �C���j �D$(P�D$P���D$H�+������L$���D$<訽����t�L$D�����"�|A�L$$���   Q�@L�ЋL$H��P�g����|A�D$$���   P�	�D$   �D$@ �ыD$H���L$4d�    Y^[��4� ����������j�h#�d�    P��(SV�8A3�P�D$4d�    ���D$    �D$$    �D$,    �D$P�L$�D$@   �D$�  �D$     �D$$    �3���j �D$(P�D$P���D$H�������L$���D$<蘼����t�L$D�����"�|A�L$$���   Q�@L�ЋL$H��P�W����|A�D$$���   P�	�D$   �D$@ �ыD$H���L$4d�    Y^[��4� ����������j�hN�d�    P��$V�8A3�P�D$,d�    ��|A�t$<�D$     �D$(    ���   �L$ �@(Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    ����j�D$ P�D$P���D$@�����L$�D$4 �z����|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�hy�d�    P��$V�8A3�P�D$,d�    ��|A�t$<�D$     �D$(    ���   �L$ �@(Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �0���j�D$ P�D$P���D$@�(����L$�D$4 蚺���|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h��d�    P��,SV�8A3�P�D$8d�    ���D$(    �D$0    �D$P�L$�D$D    �D$ �  �D$$    �D$(    �k���j �D$,P�D$P���D$L�S������L$���D$@ �й����tW��D$�D$��|A�L$(���   Q�@<�Ѓ��|A�\$�L$(���   Q� �D$D�������D$���L$8d�    Y^[��8�������������j�h��d�    P��V�8A3�P�D$$d�    ���D$4�D$   �D$�D$P�L$8�D$0    �D$�  �D$    �D$    �h���j�D$P�D$<P���D$8�`����L$4�D$, �Ҹ���|A�L$���   Q� �D$0�����Ѓ��L$$d�    Y^��(� j�h��d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     諶��j �D$$P�D$P���D$D�������L$���D$8 ������t3���|A�L$ ���   Q�@8�Ѓ����|A�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h%�d�    P��$V�8A3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    輵��j�D$ P�D$P���D$@�����L$�D$4 �&����|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�hP�d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �����j �D$$P�D$P���D$D��������L$���D$8 �`�����t:�|A�t$@���   W��	����D$ P�F�D$<�����у��K�|A�L$ ���   Q�@P���~ �t$D�|Af��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h{�d�    P��$V�8A3�P�D$,d�    ��|A�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    谳��j�D$ P�D$P���D$@�����L$�D$4 �����|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h��d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     ����j �D$$P�D$P���D$D��������L$���D$8 �P�����t:�|A�t$@���   W��	����D$ P�F�D$<�����у��K�|A�L$ ���   Q�@P���~ �t$D�|Af��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h��d�    P��$V�8A3�P�D$,d�    ��|A�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    蠱��j�D$ P�D$P���D$@�����L$�D$4 �
����|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� �������̡|A���@Lj�t$���   Q�L$Q�ЋL$$�~ f��~@f�A���� � ��̡|A���@Lj �t$���   Q�L$Q�ЋL$$�~ f��~@f�A���� � ���j�h��d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �[���j �D$$P�D$P���D$D�C������L$���D$8 �������t:�|A�t$@���   W��	����D$ P�F�D$<�����у��K�|A�L$ ���   Q�@P���~ �t$D�|Af��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h'�d�    P��$V�8A3�P�D$,d�    ��|A�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    ����j�D$ P�D$P���D$@�����L$�D$4 �z����|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�hR�d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �K���j �D$$P�D$P���D$D�3������L$���D$8 谯����t:�|A�t$@���   W��	����D$ P�F�D$<�����у��K�|A�L$ ���   Q�@P���~ �t$D�|Af��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h}�d�    P��$V�8A3�P�D$,d�    ��|A�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    � ���j�D$ P�D$P���D$@������L$�D$4 �j����|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h��d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �;���j �D$$P�D$P���D$D�#������L$���D$8 蠭����t3���|A�L$ ���   Q�@8�Ѓ����|A�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h��d�    P��$V�8A3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    �L���j�D$ P�D$P���D$@�D����L$�D$4 趬���|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�h��d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     苪��j �D$$P�D$P���D$D�s������L$���D$8 ������t:�|A�t$@���   W��	����D$ P�F�D$<�����у��K�|A�L$ ���   Q�@P���~ �t$D�|Af��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h)�d�    P��$V�8A3�P�D$,d�    ��|A�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �@���j�D$ P�D$P���D$@�8����L$�D$4 說���|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�hT�d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �{���j �D$$P�D$P���D$D�c������L$���D$8 ������t3���|A�L$ ���   Q�@8�Ѓ����|A�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h�d�    P��$V�8A3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    茧��j�D$ P�D$P���D$@�����L$�D$4 ������|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�h��d�    P��$SV�8A3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �˦��j �D$$P�D$P���D$D�������L$���D$8 �0�����t3���|A�L$ ���   Q�@8�Ѓ����|A�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h��d�    P��$V�8A3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    �ܥ��h�   �D$ P�D$P���D$@������L$�D$4 �C����|A�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� �������t��t��t3�ø   ���̡|AQ�@L�@L�Ѓ���������������̡|AQ�@L�@P�Ѓ�����������������t$�|A�t$�@L�t$���  Q�Ѓ�� ������������̡|A�t$�@LQ��  �Ѓ�� ����̡|A�t$�@LQ���   �Ѓ�� ����̡|AQ�@L�@X�Ѓ�����������������t$�|A�t$�@L�t$�@\Q�Ѓ�� j�h �d�    P��0SVW�8A3�P�D$@d�    ��|A�@L�@�Ћ؅�u�L$@d�    Y_^[��<� �L$藺���D$H    �D$(    �D$0    �D$4    �D$<    �D$8    �t$P�D$�D$0�|A�\$(�@h]  �@0�L$�D$P�С|Aj ���   j �@S���Ѕ���   �|AS�@L�@�Ћ�������   ���|A���   �΋R(�ҋ��D$$Ph�   �t$0�H�������ts�L$<��tk�|Aj ���   ���   �ЋЅ�tP�|AV���   �ʋ@<�С|A�L$<���   Q���   �Ѓ���t�|AV�@@�@�Ѓ������`����+�|AS�@@�@�С|A�L$@���   Q���   �Ѓ�3ۍL$$�D$H ������L$�D$H�����t����ËL$@d�    Y_^[��<� ������������̡|AQ�@L�@`�Ѓ���������������̡|AQ�@L�@d�Ѓ���������������̡|A�t$�@LQ�@h�Ѓ�� �������̡|AQ�@L��D  �Ѓ������������̡|AQ�@L�@l�Ѓ���������������̡|A�t$�@LQ���   �Ѓ�� ����̡|A�@L�@����̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@L���   ��Y�������������̡|AQ�@L���   �Ѓ��������������t$�|A�t$�@L�t$���   �t$�t$Q�Ѓ�� ������t$�|A�t$�@L�t$���   Q�Ѓ�� ��������������t$�|A�t$�@L�t$��   �t$Q�Ѓ�� ����������t$�|A�t$�@L�t$��   Q�Ѓ�� ������������̡|A�@L��H  ��|A�@L��L  ��|A�@L��P  ��|A�@L��T  ��|A�@L��p  ��|A�@L��t  ��|A�@L���  ��|A�@L���  ��|A�@L���  ��|A�@L���  ���T$ V�t$�D$h��hp�h`�hP�R�t$4�q�t$4�Q�t$4�|A���@L�$�t$4���   VQ�Ѓ�4^�  ����̡|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|A�@���   ��|AV�@�t$���   �6�Ѓ��    ^��������������̡|AV�@L�@�Ћ���u^á|Aj �t$�@�t$��h  �t$V�Ѓ���u�|AV�@@�@�Ѓ�3���^�������������̡|Aj �H�t$�D$�� P�t$��h  �t$�Ѓ�������̡|A�@���   ��|A�@L���   ���t$�|A�t$�@�t$���   �t$ �t$ �t$ �t$�Ѓ��j�h+�d�    P�� V�8A3�P�D$(d�    �D$    �D$    �D$    �D$    �D$    �D$$    �D$     �|A�D$0    ���   ���   �ЉD$�t$8�D$0��t<��t8�|Aj�QLP���   ���ЋD$�D$ �D$Ph=���t$�S���������   �|A�L$���   Q���   �D$4 �Ѓ��L$�D$    �D$0�����n����ƋL$(d�    Y^��,������������j�hV�d�    P�� V�8A3�P�D$(d�    �D$    �D$    �D$    �D$    �D$    �D$$    �D$     �|A�D$0    ���   ���   �ЉD$�t$8�D$0��t<��t8�|Aj�QLP���   ���ЋD$�D$ �D$Ph<���t$�3���������   �|A�L$���   Q���   �D$4 �Ѓ��L$�D$    �D$0�����N����ƋL$(d�    Y^��,�����������̡|A�@L���   ��|A�@L���   ��|A�@L��  ��|A�@L��@  ���L$�� �������̋L$�t$��P��̋L$�t$��t$�P����������������t$�L$�t$��t$�t$�P������̡|AV���   �񋀌   V�Ѓ��    ^��������������̡|AQ�@D�@$�Ѓ���������������̡|Aj �@D�t$� �Ѓ�����������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@D�@�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|A�@D� �����̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|A�t$�@Dh2  � �Ѓ��������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|Aj �@D�t$� �Ѓ�����������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|A�t$�@Dh'  � �Ѓ��������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|A�t$�@DhO  � �Ѓ��������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|A���@XQ� �L$Q�ЋL$$�~ f��~@f�A�~@f�A���� � ��̡|A���@XQ�@�L$Q�ЋL$$�~ f��~@f�A�~@f�A���� � �̡|A���@XQ�@�L$Q�ЋL$$�~ f��~@f�A�~@f�A���� � �̡|A��`�@XV�@WQ�L$Q�Ћ��D$t���   ���_^��`� �������������̡|A�t$�@XQ�@�Ѓ�� �������̡|A�t$�@XQ�@�Ѓ�� �������̡|A�t$�@XQ�@�Ѓ�� �������̡|A�t$�@XQ�@�Ѓ�� �������̡|A�t$�@XQ�@$�Ѓ�� �������̡|A�t$�@XQ�@ �Ѓ�� �������̡|Aj �@Dh�  � �Ѓ����������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@D�@(�Ѓ���������������̡|AQ�@D�@�Ѓ���������������̡|A�t$�@D�t$�@Q�Ѓ�� ���̡|Aj �@Dh:  � �Ѓ����������̡|AV�@@�t$�@�6�Ѓ��    ^�̃��|A�$    �D$    ���   �$�@Rj�����#D$��������������̡|Aj �@Dh�F � �Ѓ����������̡|AV�@@�t$�@�6�Ѓ��    ^�̋D$����u��� �D$�|A�$    ���   �$�@Rj������؃�� �̡|Aj �@Dh�_ � �Ѓ����������̡|AV�@@�t$�@�6�Ѓ��    ^�̡|AQ�@\�@�Ѓ���������������̡|AQ�@\�@�Ѓ���������������̡|A�t$�@\Q�@�Ѓ�� �������̡|A�t$�@\�t$�@Q�Ѓ�� ���̡|A�t$�@\Q�@�Ѓ�� �������̡|AQ�@\�@�Ѓ���������������̡|A�t$�@\Q�@ �Ѓ�� �������̡|A�t$�@\�t$�@$Q�Ѓ�� �����t$�|A�t$�@\�t$�@`�t$Q�Ѓ�� �����������̡|A�t$�@\Q�@0�Ѓ�� �������̡|A�t$�@\Q�@@�Ѓ�� �������̡|A�t$�@\Q�@D�Ѓ�� �������̡|A�t$�@\Q�@H�Ѓ�� �������̡|AQ�@\�@4�Ѓ���������������̡|A�t$�@\�t$�@8Q�Ѓ�� ���̡|A�t$�@\Q�@<�Ѓ�� ��������QSUVW�|$��j ���|����|AU�@\�@�Ѓ���S���a���3���~G�	��$    ���|A�L$�@\Q�@`�L$Qh���VU�Ѓ����t$�$����t$������F;�|�_^][Y� �����������̃�S�\$W�D$��P�������|$ ��   �|AW�@\�@�Ѓ��D$P�������D$��taV3���~L���D$P���Ԩ���D$P���Ȩ���L$;L$!�|AQ�@\W�@�ЋL$$A���L$;L$~�F;t$|�^_�   [��� _�   [��� ����������̡|A�@\� �����̡|AV�@\�t$�@�6�Ѓ��    ^���    �A    �A    �A    �����V��V�u���FP�~u�����F    �F    ^������������S�\$V��W�~�    �    �F    �F    �CV;C��   �(u��W�"u���F    �F    �|Ah�	�@jI���   j�Ѓ������   �|Ah�	�@jN���   j�Ѓ����uV��t������_^[� ��F   �F   ����C�A��C�A�_�    ��^[� �t��W�|t���F    �F    �|Ah�	�@jI���   j�Ѓ����tZ�|Ah�	�@jN���   j�Ѓ�����Z�����F   �F   ����C�A��C�A��C�A��    _��^[� ����������V�t$���    �F    �F    �F    �  ��^� ���V�t$���  ��^� ��������������SUV��V�s���nU�|s���\$���F    �F    ��t(�|Ah�	�H��    jIP���   �Ѓ����u^]3�[� W�|$��t;�|Ah�	�H��    jNP���   �Ѓ��E ��uV��r����3�_^][� �~_�^^]�   [� �������������V��V��r���FP�r�����F    �F    ^������������SV��WV�r���^S�r���|$���F    �F    ����   �? ��   �W����   �|Ah(
�H��    jlP���  �Ѓ����t<� t>�W��t7�|AhT
�H��    jqP���  �Ѓ����u���'���_^3�[� �G�F�G�F��P�7�6��'  �����t�F��P�wQ��'  ��_^�   [� ���������������SUV��WV�q���~W�q�����|$ �F    �F    ��   �\$����   �|Ah�
�@��    ���  h�   Q�Ѓ����tB�l$ ��tL�T$��tD�|Ah�
�H��    h�   P���  �Ѓ����u���&���_^]3�[� �D$�F�,�F   �|Ah�
�@h�   ���  j�Ѓ����t���    P�t$ �^�6�&  ����t�F��PU�7�&  ���   _^][� ��_^]�   [� ��������������    �A    �A    �A    �����U������   �U��V�HWW�3��<��D$�|$@�L$}
��_^��]� ����  �0�U�f(ύ@�F�~ʍ@f(��D��,��t��\D��D$�\t��8�L$(�|$ �T$�\$0�\��D$8����   ��������f(ƍ@f(��$��T��\T��\��\��\\����Y��Y��Y��Y��\�f(��Y��Y��XL$(�\�f��\$0�\��L$(�Xl$�Xt$ �l$f�f(��D$ f�O�f����T$W��(��YL$(�YD$ �}f�?�X�f(��Y�f�f��X���$  �T$(�\$ f(�W�f.͟��Dz�L$f(�f(�f(��&���^��L$f(�f(��Y��Y��Y�f�gH�%�	fT�fT�f/�f�wPf�GX��   f(�fT�f/���   �GH�WX�gP(��Y�(��Y��\��Y��\�f�_�\�f�O f�g(�OX�P�Y(�W�gH(��YG (��YWP�\�(��YG(�Yg �Y�f�0�\��\�f�_8f�g@�)  �WPfT�f/��_X��   �OH�Y�f(��Y��\��\��Y�f�Gf�_ �\�f�O(�(�G �YGX�YP�O�wH(��Y_X�YOP�\�f(��YG(�Yw f�0�\��\�f�_8f�w@�   f(��Y�(��Y��\��GH�Y�f�O0�\��\�f�_8f�G@�oP�X�Y8�OH�w0(��YG@(��Y_@�YO8�\�(��YGX�Y�f��\��\�f�_ f�w(�D$`WP����U���D$�   ���W�3�3Ʌ�~w��r]�p��W�W�%  �yH���@��+���    �o���f���oD��f��;�|�f��fo�fs�f��fo�fs�f��f~ϋt$;�}�F<�A;�|���t$�M��u�A0�D$(���q �@�D$    ���d��\��Y�f(��YI�D$(�Y��X	�D��Xq�@�X��AH�Y��X��A8�Y��L$ �I(�X��AP�Y��Y��T��X��A@�XI�Y��$��X��AX�Y�(��YY�X�(��YA0�Xf�L$X�L��D$�X�(��YAH�@���X�(��YA8�YQ@�\$(��YY �Ya(�D$�XY�Xa�X�(��YAP�YIX�X��X��X��\$0f�d$8���  3�������|$�D$(׋��@�,��T��L�f(��Ya(��YA0�X!f(��YY �Yi(�X��XY(��YAH�Xi�D$@�X�(��YA8�YQ@�D$�X�(��YAP�YIX�X��T$0�X�(��X�f(��\��\��\�f�\$0�YL$�YD$ �Y��X��~D$�D$ �~D$8f�D$X�X�f�f�d$f�l$8�X�;D$������|$@�D$@_^��]� �����������̋�����������T$�   @t������@��wm�$���D$� ����D$� ���� �
�D$��D$�J�� �J�D$��D$�J�� �J�D$��D$�J�� �J�D$��D$�
�� �I ����˵���S��V�����%���W��   @t�����ʃ��|$;�t�����t�t$�����t��t$;�t>�����t6�΁����Eǃ��t����   �_�^�[� ��   ���Ё�   @�_^[� ���U�������AW�SVf(�f(�f(�W�L$�\$�T$ �D$���L  �9�u������Ш�)  ���������U��Z�@�[�<��l��\<��\l�;Zuc�\��B�\\��@�d��\d��T��\T��4��\4�f(��Y�f(��Y��Y��\�f(��Y��\��Xd$(��d�d��B�\d��@�B�@�T��\��\\��\T��4��\4�f(�f(��Y��Y��Y��\�f(��Y��\��X\$�XL$�Y��Y��\$�L$�\��Xt$ (��T$ ���L$�����f(��Y�f(��Y��X�f(��Y��X��  f(�W�f.П��D�Ez� �@�@_^[��]� ���^�_^[(��YD$� (��YD$�@�D$�Y��@��]� ���������U������<���5��AS3�Vf�f�f�f�W�D$�L$�|$ �t$(�l$0�d$8�T$@�D$���4  ��u��    ������Ш��  ���������M��@��ts��f/�v
f(��D$�\�f/�v
f(��L$�\�f/�v
f(��|$ f/�v
f(��t$(�T�f/�v
f(��l$0f/�vPf(��D�~4��~l��~d�f�f�f�   �t$(�l$0�D$�L$�|$ �T$@�d$8�A�@��ts��f/�v
f(��D$�\�f/�v
f(��L$�\�f/�v
f(��|$ f/�v
f(��t$(�T�f/�v
f(��l$0f/�vPf(��D�~4��~l��~d�f�f�f�   �t$(�l$0�D$�L$�|$ �T$@�d$8�y���ts��f/�v
f(��D$�\�f/�v
f(��L$�\�f/�v
f(��|$ f/�v
f(��t$(�T�f/�v
f(��l$0f/�vPf(��D�~4��~l��~d�f�f�f�   �t$(�l$0�D$�L$�|$ �T$@�d$8�A;�t8�@�L$��P�E  �T$@�d$8�l$0�t$(�|$ �L$�D$���L$�@�����te�Ef(��X�f(��X��P	f(��X��Y��Y��Y�f�f�Pf�H�\0�\h�\`�Ef�0f�hf�`_^[��]� �EW�f� f�@f�@�E_f� ^f�@f�@[��]� ��������̋Q3���|�	��t��~�    t@��Ju��3����������̋QV�t$��;�}�	���    u@��;�|����^� +�@^� ���������������VW�|$���x*���t$�v3Ʌ�~��I ���%���;�tA��;�|�_���^� _��^� �����������SV�q2ۅ�~;�W�|$�
����%���;�u��   @u�����t	�   ���3�
؃�Nu�_��^��[� V�q3҅�~�	�d$ ��   @u	�����tB��Nu��^�����V�q3҅�~�	�d$ ����ШtB��Nu��^�����������QV��3�9N~��I �A�d�����;N|��N��~gSU3�W�   �T$����x;���������;�},�I ����<����������;�u��   ��@;F|ۋT$�NE���E��T$;�|�_][^Y����������������h�Ajh_� �  ����uË@����V�t$�> t1h�Ajh_� �  ����t��L$�@�L$Q�Ѓ��    ^����Vh�Ajh_� ���\  ����t�@��t�t$����^� 3�^� ������������Vh�Ajh_� ���  ����t�@��t�t$����^� 3�^� ������������Vh�Ajh_� ����  ����t�@��t�t$���t$�t$��^� 3�^� ����Vh�Ajh_� ���  ����t�@��t�t$����^� 3�^� ������������Vh�Aj h_� ���\  ����t�@ ��t�t$����^� 3�^� ������������Vh�Aj$h_� ���  ����t�@$��t�t$����^� 2�^� ������������Vh�Aj(h_� ����  ����t�@(��t��^��3�^������Vh�Aj,h_� ���  ����t�@,��t��^��3�^������Vh�Aj0h_� ���|  ����t�@0��t�t$����^� 3�^� ������������Vh�Aj4h_� ���<  ����t�@4��t�t$���t$��^� ���^� �������Vh�Aj8h_� ����  ����t�@8��t��^��3�^������Vh�Aj<h_� ����  ����t�@<��t�t$����^� ��Vh�Aj@h_� ���  ����t�@@��t�t$����^� ��Vh�AjDh_� ���l  ����t�@D��t�t$����^� 3�^� ������������Vh�AjHh_� ���,  ����t�@H��t�t$����^� ��Vh�AjLh_� ����  ����t�@L��t��^��3�^������Vh�AjPh_� ����  ����t�@P��t��^��3�^������Vh�AjTh_� ���  ����t�@T��t��^��^��������Vh�AjXh_� ���l  ����t�@X��t��^��^��������Vh�Aj\h_� ���<  ����t�@\��t��^��^��������Vh�Aj`h_� ���  ����t�@`��t�t$���t$��^� 3�^� ��������Vh�Ajdh_� ����  ����t�@d��t�t$���t$��^� 3�^� ��������Vh�Ajhh_� ���  ����t�@h��t�t$���t$�t$�t$�t$��^� ��Vh�Ajlh_� ���L  ����t�@l��t�t$���t$�t$��^� 3�^� ����Vh�Ajph_� ���  ����t�@p��t�t$���t$��^� 3�^� ��������Vh�Ajth_� ����
  ����t�@t��t�t$���t$��^� 3�^� ��������Vh�Ajxh_� ���
  ����t�@x��t�t$���t$��^� 3�^� ��������Vh�Aj|h_� ���L
  ����t�@|��t�t$����^� 3�^� ������������Vh�Ah�   h_� ���	
  ����t���   ��t�t$���t$��^� 3�^� ��Vh�Ah�   h_� ����	  ����t*���   ��t �t$���t$�t$�t$�t$�t$��^� ���^� �Vh�Ah�   h_� ���y	  ����t*���   ��t �t$���t$�t$�t$�t$�t$��^� ���^� �Vh�Ah�   h_� ���)	  ����t"���   ��t�t$���t$�t$�t$��^� 3�^� ����������Vh�Ah�   h_� ����  ����t���   ��t�t$����^� 3�^� ������Vh�Ah�   h_� ���  ����t���   ��t�t$����^� ������������Vh�Ah�   h_� ���Y  ����t���   ��t�t$���t$��^� 3�^� ��Vh�Ah�   h_� ���  ����t���   ��t�t$���t$�t$��^� 3�^� �������������̃��L$�T$�D$�R�X�A�\B�\��\Y�Y �Y�Y�X��X��$�$�������h�A�t$h_� �}  �����������̃y0 �D$tq��f/�v�	�H�Af/�v�I�H�Af/�v�I� f/Av�A�@f/A v�A �@f/A(vI�A(� �~ f�A�~@f�A �~@f�A(�~Af��~A f�A�~A(f�A�A0   � ̡|A�@d�@P����̋L$�9 t�|A�L$�@d�@T���������t$�|A�t$�@h�t$� �t$Q�Ѓ�� ��������������t$�|A�t$�@h�t$���   �t$Q�Ѓ�� ����������t$�|A�t$�@h�t$�@Q�Ѓ�� �t$�|A�t$�@h�t$�@ �t$�t$Q�Ѓ�� ���������t$�|A�D$�@h�����   �$Q�Ѓ�� ��������t$�|A�D$�@h�����   �$Q�Ѓ�� ������̡|A�t$�@h�t$���   Q�Ѓ�� ̡|A�t$�@h�t$���   Q�Ѓ�� ��D$�|A���@h�t$<���   �t$<���D$�D$@�$�t$<�t$<Q�L$$Q�ЋL$D�~ f��~@f�A�~@f�A����@�$ ������D$�|A���@h�t$8���   ���D$�D$<�$�t$8�t$8Q�L$ Q�ЋL$@�~ f��~@f�A�~@f�A����<�  ���������j�h��d�    P��VW�8A3�P�D$$d�    ���D$    �|$4�    �G    �D$8�D$�D$P�L$�D$0    �D$   �D$     �D$$    �Jm��j W�D$P���D$8   �3����L$�D$, �n���ǋL$$d�    Y_^��$� ����������������t$�|A�t$�@h�t$���   �t$Q�Ѓ�� ��������̡|A�t$�@hQ���   �Ѓ�� ����̡|A�@h�@X����̋L$�9 t�|A�L$�@h�@\�������̡|A�@h���   ��|A�@h���   ��|A�@h���   ���t$�|A�t$�@h�t$�@`�t$�t$�t$�t$Q�Ѓ� � �t$�|A�t$�@h�t$�@d�t$�t$�t$�t$Q�Ѓ� � �|A�t$�@h�t$�@hQ�Ѓ�� ���̡|A�t$�@h�t$�@lQ�Ѓ�� ���̡|A�t$�@h�t$�@pQ�Ѓ�� �����t$�|A�t$�@h�t$���   �t$�t$�t$�t$Q�Ѓ� � ��������������t$�|A�t$�@h�t$���   �t$�t$�t$�t$Q�Ѓ� � ��������������t$�|A�t$�@h�t$���   �t$�t$�t$�t$Q�Ѓ� � ��������������t$�|A�t$�@h�t$���   �t$�t$Q�Ѓ�� ������t$�|A�t$�@h�t$���   �t$Q�Ѓ�� ����������t$�|A�t$�@h�t$�@tQ�Ѓ�� �|A�t$�@hQ�@x�Ѓ�� �������̡|A�@h���   ���t$�|A�t$�@h�t$�@|Q�Ѓ�� �t$�D$�|A���@h�D$�D$(���   �D$�D$ �$Q�Ѓ� � ��������������̋L$�D$Q��D$j�t$�A胎�������������������̸   �����������V�t$��t���u7j�t$�f�������u3�^Ë������ȅ�t��t��D$3�;AOʋ�^�;8Au���T  ��%� U���EV��t%Wh���~��7jV�'  �EtW�7@��Y��_���  �EtV� @��Y��^]� ��������Vh�   �< Y��V� ��D��D��u3�@^Ã& �  h��D  �$8��8  Y3�^�U��QQ�} SVW�)  ��A���  H��Ad�   3��P�}���D�;�t3�������u���E�   �=�Dtj�  Y�  �5�D� ���u����   �5�D� �؉u�]��;�r\9;t�W� 9t��3� W��� ����5�D�5 ���5�D�E��֋M�9Mu�u9Et���M�u�E��띃��tV�� YW� ��D��D��D�=�D9}���   3���   3��   �}��   d�   3��P����D�;�t3�������u��3�F9=�Dj_t	j�  �5h� h� ��D   �  YY��u�h� h� �   Y�=�DY��u3���=�D th�D�  Y��t�uW�u��D��A3�@_^[�� U��}u��  �u�u�u�   ��]� jh.�  3�@���u�3ۉ]��}�=@A�E���u9=�A��   ;�t��u8���t�uW�u�Ћ��u����   �uW�u�������u����   �uW�u�:|�����u��u.��u*�uS�u� |���uS�u�@������t	�uS�u�Ѕ�t��uK�uW�u�������#��u�t4���t+�uW�u�Ћ���M�� �E�QP�c  YYËe�3ۋ�u�]��E������   ����  Ëu��@A�������%� �=�D t3��Vjj �P YY��V� ��D��D��ujX^Ã& 3�^�jh0.�:  �5�D�5 �։E���u�u�X Y�ej�  Y�e� �5�D�։E��5�D�։E��E�P�E�P�u�5 ��P�e  �����}��u��֣�D�u��֣�D�E������   ����  Ë}�j�%  Y�U���u�P��������YH]��%� �%| �%x �%L �%$ �%( �%, U��� j��D��  �u��  �=�D YYuj��  Yh	 ���  Y]�U���$  j��  ��tjY�)��B��B��B��B�5�B�=�Bf��Bf��Bf��Bf��Bf�%�Bf�-|B���B�E ��B�E��B�E��B��������A  ��B��A��A	 ���A   ��A   jXk� ǀ�A   jXk� �8A�L�jX�� �<A�L�h�������jhP.�   �e� �]�Ë}�ǋu��u�e� O�}x+�u���U��3�@�E��E������   �!  � �}�]�u�E��u�uWSV�   �jhp.�  �e� �Mx:�M+M�M�U��E�E�E� �E��E��8csm�t�E�    �E���  �e��E������  � ��%0 �%4 �%8 ������������U��ES�H<�V�A�Y��3��W��t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�h�.h��d�    P��SVW�8A1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��E�MZ  f9t3�]ËH<�3��9PE  u�  f9Q��]�U����8A�e� �e� VW�N�@��  ��;�t��t	�У<A�f�E�P� �E�3E�E��  1E�� 1E��E�P� �M�3M�E�3M�3�;�u�O�@����u��G  ��ȉ8A�щ<A_^��VW��������t�Ѓ�;�r�_^�VW� � ����t�Ѓ�;�r�_^���%@ �%D h�D�   Y�������������h��d�5    �D$�l$�l$+�SVW�8A1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�U���u�u�u�uh��h8A�5   ��]��%H �%� �%T �%` �%d �%h �%l �%p �%t �% �������̍M��88���M�頋���M��(8���T$�B؋J�3������������������������h�jEh�A�E�P��7����ËT$�B��J�3��N�����T��������������̍M��7���M��P]���M��H]���M��7���T$�B��J�3������T��������̍M��x7���M��p7���T$�B؋J�3�����������������̍M���\���T$�B��J�3������d����hj;h�A�E�P�(7����ËT$�B��J�3��{����@�����M���6���M���6���EЃ��   �e���M��6��ËT$�BЋJ�3��7�����=����M��6���M��6���EЃ��   �e���M�6��ÍM��6���T$�BЋJ�3��������������M��a6���M��Y6���EЃ��   �e���M�A6��ÍM��86���M��06���T$�BЋJ�3������������M��6���M��6���EЃ��   �e���M��5��ÍM���5���M���5���M���5���T$�BЋJ�3��;������A����M��5���E����   �e���M��5��ËE����   �e���M��5��ËT$�B��J�3��������������M��\5���E����   �e���M��D5��ËE����   �e���M��+5��ËT$�B��J�3������h������������������̍M���4���E����   �e���M��4��ËT$�B�J�3��F������L������̍M��XZ���Eԃ�t�e���M�DZ��ËT$�B��J�3��
����$�����������̋M��x4���T$�B��J�3��������������M��U4���T$�B��J�3�������������M��24���T$�B��J�3������������M��4���T$�B��J�3��v������|����M���3���T$�B��J�3��S����h�Y����M���3���E����   �e���M�3��ËT$�B�J�3������D�����M��-Y���M�3���Eԃ��   �e���M�Y��ÍM��d3���T$�B؋J�3������� ������M���X���M�93���Eԃ��   �e���M��X��ÍM��3���T$�B؋J�3������������M��X���Eԃ��   �e���M��2��ÍM���2���T$�B��J�3��;������A����M�2���E����   �e���M�9X��ËT$�B��J�3�������������M��u2���E����   �e���M�]2��ËT$�B�J�3��������������M��92���T$�B�J�3������l�����M��2���T$�B�J�3��}����H�����M���1���T$�B�J�3��Z����$�`����M��pW���M��1���Eԃ��   �e���M�PW��ÍM��1���T$�B؋J�3������ �����M��$W���M�|1���Eԃ��   �e���M�W��ÍM��[1���T$�B؋J�3��������������M��81���E����   �e���M� 1��ËT$�B�J�3������������M��V���M���0���T$�B��J�3��[������a����M��qV���M��0���Eԃ��   �e���M�QV��ÍM��0���T$�B؋J�3������p�����M��%V���M�}0���Eԃ��   �e���M�V��ÍM��\0���T$�B؋J�3�������L������E����   �e���M���U��ÍM�� 0���E����   �e���M��U��ËM��/���E����   �e���M�U��ÍM���/���M���/���T$�B��J�3��=����(�C����M��SU���M�/���Eԃ��   �e���M�3U��ÍM��/���T$�B؋J�3�������������M��g/���E����   �e���M�O/��ËT$�B�J�3�������������̍�h�����T����X����/���M��T���M��T���M��T���M��T���T$��\�����X���3��[����T�a�����������̍M���.���E����   �e���M�.��ËT$�B�J�3������������M��<����T$�B�J�3��������������M������E����   �e���M����ËT$�B�J�3������������M����ʖ���T$�B��J�3������d����hPh�   h�A�E�P�.����ËT$�B��J�3��Z����@�`����M���m����T$�B��J�3��4�����:����M��*k���M��-���T$�BЋJ�3��	���������������̍M���j���T$�BЋJ�3�������P!������M���j���T$�B�J�3������,!������E����   �e���M�ҕ��ÍM��ɕ���T$�B�J�3������!�����M��vj���M�鞕���T$�BԋJ�3��U����� �[����M��Kj���M��s����T$�B��J�3��*����� �0����M�� j���M��H����T$�B��J�3�������� �����M���i���M������T$�B؋J�3�������x ������M��J,���T$�B�J�3������T �����M��',���T$�B�J�3������0 �����M��,���M���+���T$�B܋J�3��c���� �i����M��yQ���M��qQ���M���+���T$�B��J�3��0������6����M��+���T$�B�J�3������������M��#Q���T$�B��J�3��������������M���h���M������M�� ����M�������T$�B؋J�3������|�����M��h���T$�B�J�3������X�����M��h���T$�B�J�3��i����4�o����M��_h���T$�B�J�3��F�����L����M��<h���M��d����T$�B؋J�3��������!����M��h���M��9����T$�B؋J�3��������������M�������T$�B��J�3��������������M��C*���T$�B��J�3������������M�� *���T$�B��J�3������\�����M���)���T$�B�J�3��d����8�j����M���)���T$�B�J�3��A�����G����M��)���E����   �e���M�)��ËT$�B�J�3������������EЃ��   �e���M�k)��ÍM��b)���M��Z)���T$�BȋJ�3��������������M��7)���M��/)���M��')���M��)���M��f���M��)���T$�B��J�3��v������|����M���(���T$�B��J�3��S������Y����M���(���M���(���M��(���M��1f���T$�B��J�3������`�����M��f���M��f���T$�B��J�3�������<������M���e���T$�B�J�3�������������M��@(���M��8(���M��0(���T$�BȋJ�3������������M��(���T$�B��J�3��t������z����̋M���镐���M�鍐���T$�B�J�3��D����"�J����̋E����   �e���M�'��ËT$�B��J�3����������������������̍M�x'���T$�B��J�3�������H"�����������������̍M���d���E܃��   �e���M�d��ËT$�B�J�3�������!�������̍M��L���Eԃ��   �e���M�L��ËT$�B��J�3��V�����!�\������̍M��Hd���T$�B�J�3��/����t"�5���������������̍M���N���E���   �e���M�N��ËT$�B��J�3�������D#������M��N���E���   �e���M�tN��ËT$�B��J�3������ #�����M��PN���E܃��   �e���M�8N��ËT$�B�J�3��n�����"�t����E����   �e���M��%��ÍM���%���T$�B�J�3��2�����"�8����M�HK���T$�B��J�3������p#����������������̋E���t�e���M�l%��ËT$�B��J�3�������T'������M��H%���M��@%���T$�B��J�3������0'�����M��%���E����   �e���M�%��ËT$�B�J�3��k����'�q����M���$���E����   �e���M��$��ËT$�B�J�3��/�����&�5����E���t�e���M�9J��ËT$�B��J�3��������&�����E���t�e���M��a��ËT$�B��J�3��������&������M��E$���E����   �e���M�-$��ËT$�B�J�3������|&�����M��	$���E����   �e���M��#��ËT$�B�J�3��W����X&�]����M��mI���Eԃ�t�e���M�#��ËT$�B��J�3������4&�%����M��E����E����   �e���M�-���ËT$�B�J�3�������&������M���`���M������Ẽ��   �e���M�`��ËT$�BԋJ�3�������%�����M��#���E����   �e���M��"��ËT$�B�J�3��c�����%�i����M�鉋���E����   �e���M�q���ËT$�B�J�3��'�����%�-����M��`���T$�B܋J�3�������%�
����Ẽ��   �e���M�j"��ÍM���_���M��	����T$�BЋJ�3�������\%������Ẽ��   �e���M�&"��ÍM��_���M��Ŋ���T$�BЋJ�3��|����8%�����M��r_���M�隊���T$�B؋J�3��Q����%�W����M��G_���M��o����T$�B؋J�3��&�����$�,����M��_���E܃�t�e���M�_��ËT$�B�J�3��������$����������������̍M���^���E܃�t�e���M��^��ËT$�B�J�3�������-�����M��^���E܃�t�e���M�^��ËT$�B�J�3��r�����-�x����M�阉���M��I���T$�BԋJ�3��G����h-�M����M��m����M���H���T$�B؋J�3������D-�"����M��B����M��H���Ẽ��   �e���M�F��ËT$�BЋJ�3������� -������M�������M��vH���Ẽ��   �e���M��E��ËT$�BЋJ�3�������,�����M�麈���M��2H���T$�B؋J�3��i�����,�o����M�鏈���M��H���T$�B؋J�3��>�����,�D����M��d����M���G���T$�B̋J�3�������,�����M��9����M�G���T$�B��J�3�������l,������M������M��G���T$�BԋJ�3������H,������M������M��[G���T$�B؋J�3������$,�����M�鸇���M��0G���T$�BԋJ�3��g���� ,�m����M�鍇���M��G���T$�B؋J�3��<�����+�B����M��b����M���F���T$�BԋJ�3�������+�����M��7����M��F���T$�B؋J�3��������+������M������M��F���T$�BԋJ�3������p+������M������M��YF���T$�B؋J�3������L+�����M�鶆���M��.F���T$�BԋJ�3��e����(+�k����M�鋆���M��F���T$�B؋J�3��:����+�@����M��`����M���E���T$�BԋJ�3�������*�����M��5����M��E���T$�B؋J�3��������*������M��
����M��E���T$�BԋJ�3�������*�����M��߅���M��WE���T$�B؋J�3������t*�����M�鴅���M��,E���T$�BԋJ�3��c����P*�i����M�鉅���M��E���T$�B؋J�3��8����,*�>����M��^����M���D���T$�BԋJ�3������*�����M��3����M��D���T$�B؋J�3��������)������M���Y���M��@[���T$�BċJ�3�������)�����M��[���M�酧���T$�B܋J�3�������)�����M���Z���M��Z����T$�B܋J�3��a����x)�g�����������������̋E܃��   �e���M�h���ÍM���C���T$�B��J�3�������-��������h�������Y����̃=XA uK�PA��t�|AQ�@<�@�Ѓ��PA    V�5\A��t����@��V�'�����\A    ^�                                                                                                                                                                                                                           �1 �1 �1 �1 �1 �1 z1 2     �/ 0  0 :0 R0 d0 r0 �0 �0 �0 �/ �0 �0 �0 �0 �0 �0 1 (1 <1 `1 �/ �/ �/ �/ �/ �/ �0 �/         ��        0���            �������N���������������C-DT�!	@-DT�!�?Ocontainer.png  Ocontainer  �������N    ���������������C-DT�!	@-DT�!�?p � ` � 0 �  @b Pb `b pb �b �b �b �b �b �b P(`(�) *�+�/�/�/�/�/�/�/ 00 000src/ContainerObject.cpp 333333�?ffffff�?      �?     �o@../../resource/_api/c4d_resource.cpp    ../../resource/_api/c4d_resource.cpp    #   #   #   #   #   #   #   #   #   #   M_EDITOR    M_EDITOR    \�5 ../../resource/_api/c4d_file.cpp    ../../resource/_api/c4d_file.cpp    �������N���������������C-DT�!	@-DT�!�?res �������N    ���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  �������N���������������C-DT�!	@-DT�!�?p:\applications\maxon\cinema 4d r14.041\resource\_api\c4d_misc/datastructures/basearray.h       ~   Progress Thread 0%  ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp %   ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp �������N    ���������������C-DT�!	@-DT�!�?�� 0| @| P| `| p| �| �| �|  } } ��  � �  � 0� @� P� `� p� L�  � �  � 0� @� P� `�  � p�  � �  � 0� @� P� `� � ��  � �  � 0� @� P� `� p� �� �� ��  � �  � 0� @� `� p� �� �� -DT�!	@      Y@     �f@     @�@��������������������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  �p`    ����MbP?�������N���������������C-DT�!	@-DT�!�?        �������?-DT�!�?      �-DT�!��               �       �../../resource/_api/c4d_pmain.cpp   ../../resource/_api/c4d_pmain.cpp   %s     p:\applications\maxon\cinema 4d r14.041\resource\_api\c4d_general.h ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp              �?   ����A  4&�kC �Ngm��C  4&�k�        ��������������0�t�t����    �������N���������������C-DT�!	@-DT�!�?../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   x��    �A�AH                                                           8A��              p|�     @       ����    @   `@        ����    @   �           ��               ��|�    0@       ����    @   �            L@           ,@�|�    L@       ����    @               @�            l@�           ���    l@       ����    @   ��@        ����    @   �           ��                �@�            �@           (0    �@        ����    @               �@`           p|�    �@       ����    @   `            �@�           ����    �@       ����    @   �            �@�               �@        ����    @   �            AD           T\    A        ����    @   D             A�           ��     A        ����    @   ��� (� i� �� �� � <� �� ��  � |� �� &� q� �� �� �� � A� d� �� �� 8� |� �� �� � :� ]� �� �� 1� \� �� �� z� �� � V� �� ��  � &� ]� �� �� �� �� 7� b� �� �� �� � )� T� �� �� �� � +� N� q� �� �� �� � 0� S� v� �� �� A� d� �� �� ��  � C� s� �� �� !� a� �� �� � I� �� �� �� � L� �� �� �� $� `� �� �� � T� �� �� �� ;� f� �� �� � E� p� �� �� #� N� y� �� �� �� %� P� {� �� �� �� '� R� }� �� �� �� )� T� � �� ��  � +� V� ��                     ����P�"�                          ������    ��    ��������"�   4                       ������������"�   x                       �����    ������    �"�   �                       ����#����� �������������   �������������   ������g�    W�   _�������    ��   ��   ��"�                           "�                          "�   �                       "�   �                       "�   H                       "�   0                       "�   �                       "�   �                       ������    ��   ��   �   �����K�    ;�   C�   d�   l�   t�����X�    P�"�   �                       ������    ��"�                          ����U�����2����������\�����9������������������������    ������L�����T������    �������    ��������    ��������    �����[�    S�    t�������    ��   ��    ��������    ��   ��    ��������    w�   �    ��������    ��   ��    ��������    x�   ��    �������    �   �    0�������    ��   ��    ��"�   �                       "�                           "�                          "�                           "�   @                       "�   �                       "�   �                       "�   `                       "�   �                       "�   H                       "�   P                       "�   X                       "�   �                       "�   �                       "�   �                       "�   �                       "�   �                       "�   �                       "�   `                       "�   h                       "�   p                       "�   x                       "�   �                       ����Q�    �   (�   0�   I�   j�    r�"�   x                       ���� �    +�   6�   >�   F�   N�����x�����A������������������������������    ��������    ��"�   �                       "�   �                       "�   �                       "�   �                       "�   �                       "�   �                       "�   �                       ������"�   �                       ����;�����������\�����n�����K�����(����������������i�����F�����#�����������������!�������������������������������������    ��������    ��������    ������D�    L�������    ��������    ������}�    ������R�    Z������    /������    �   �������    ��    ������o�    w�   ������    ��   ��������������    ��    ��     �"�                           "�   H                       "�   (                       "�   �                       "�   �                       "�   0                       "�   t!                       "�   `                       "�   �                       "�   8                       "�   @                       "�   H                       "�   P                       "�   X                       "�   �                       "�   �                       "�   `                       "�   h                       "�   p                       "�   �                       "�   x                       "�   �                       "�   x                       "�   �                       "�   �                       "�   �                       "�   �                       "�                          "�                          "�   (                       "�   8                       "�   �                       "�   �                       ��������������!�����)�����1�   9�����H�    @�"�   �!                       �����     �"�   �!                       ����`�    k�"�   "                       ������"�   @"                       ������"�   l"                       ����d�    }�����0�    (�������    ��������    ��"�   �"                       "�   �"                       "�   �"                       "�   �"                       ������"�   h#                       ������������������������������    ��������    ������V�    ^�����w�    o�����;�    3�������    ��������    {�����G�    ?������    �����o�    g�����3�    +������    +�   3�������    ��   ������ �    ������������    ��   ��    ��"�   �#                       "�   �#                       "�   �#                       "�   d$                       "�   |$                       "�   �#                       "�   �#                       "�   �#                       "�   �$                       "�   $                       "�   $                       "�   $$                       "�   4$                       "�   �#                       "�   �#                       "�   D$                       "�   T$                       "�   �$                       "�   �#                       ����F�    N������    #�������    ��������    ��������    ������o�    w�����D�    L������    !�������    ��������    ��������    ������m�    u�����B�    J������    �������    ��������    ��������    ������k�    s�����@�    H������    �������    ��������    ��������    ������i�    q�����>�    F�������    ������`�    h�����0�    (�������    ������
�    ��   �������    ��   ��"�   x'                       "�   �'                       "�   �'                       "�   �'                       "�   �'                       "�   �'                       "�   �'                       "�   �'                       "�   �'                       "�   (                       "�   (                       "�   ((                       "�   8(                       "�   H(                       "�   X(                       "�   h(                       "�   x(                       "�   �(                       "�   �(                       "�   �(                       "�   �(                       "�   �(                       "�   �(                       "�   �(                       "�   �(                       "�   H)                       "�   `)                       "�   )                       "�   )                       "�   ()                       "�   8)                       ������    ��"�   �-                       ����    ����    ����    ��    ��������    ����    ����    ��    ����    ����    ����    w�    ����    ����    ��������    ����    ����    ��������/         ,0 $  �.         *2                        �1 �1 �1 �1 �1 �1 z1 2     �/ 0  0 :0 R0 d0 r0 �0 �0 �0 �/ �0 �0 �0 �0 �0 �0 1 (1 <1 `1 �/ �/ �/ �/ �/ �/ �0 �/     x__CxxFrameHandler3  �free  malloc  ,memset  �floor (memcpy  k_libm_sse2_asin_precise m_libm_sse2_cos_precise  s_libm_sse2_sqrt_precise Q_CIfmod 1_purecall MSVCR110.dll  p ??1type_info@@UAE@XZ  s__CppXcptFilter _amsg_exit  �_malloc_crt �_initterm �_initterm_e |_lock �_unlock +_calloc_crt �__dllonexit "_onexit 
_vsnprintf  K_crt_debugger_hook  �__crtUnhandledException �__crtTerminateProcess ;?terminate@@YAXXZ �__clean_type_info_names_internal  p_except_handler4_common <EncodePointer DecodePointer �IsDebuggerPresent �IsProcessorFeaturePresent <QueryPerformanceCounter $GetCurrentProcessId (GetCurrentThreadId  �GetSystemTimeAsFileTime KERNEL32.dll              ���Q    r2          h2 l2 p2 @N �2   containerobject.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                      .?AVNodeData@@      .?AVBaseData@@      .?AVObjectData@@        .?AVContainerObject@@       .?AVSubDialog@@     .?AVGeDialog@@      .?AVGeUserArea@@        .?AVGeModalDialog@@     .?AViCustomGui@@        .?AVNeighbor@@      .?AVC4DThread@@     .?AVtype_info@@ N�@���D����                                                                                                                                                                                               �   -0s0�0131C1U1g1z1�1�1�1�1�12Q2�2�2�2�2�3�3�3�3�3 4C4T4r4�4�4�4s5�5�56/6Y6|6�6�6(7 8$8(8,8084888<8@88�89!9K9�9�9:H:j:�:;);�;�;�; <<6<g<�<�=�=>:>P>U>y>�>�>�>?!?F?u?�?�?       0c0q0�0�0;1c1�1�122C2T2o2y2�2�2�2�2�2�2�2383R3�3�3�3�34$4?4I4U4h44�4�4�4�4�45"5g5�5�5�5�5�5�56<6N6b6�6�6�6�6�6�67"7<7O7Z7~7�7�7�78&898D8h8�8�8�8�8�8�8 9:9\9y9�9�9�9�9::%:8:O:b:|:�:�:�:�:�:7;T;f;y;�;�;�;�;<<1<<<`<z<�<�<�<�<�<='=I=f=x=�=�=�=T>i>�>�>�>�>?"?*?A?�?�?   0  0  0N0w0�0�011*121I1�1�12P2y2�2�23"3+343F3Q3k3�3�3�3�3�3�324B4a4q4�4�4�455!515A5Q5a5q5�5�5�5�5�5�566)676s6�6�6�6�6�677'7=7s7�7�7�7�7�788/8a8�8�8�8�8�8�899a9�9�9�9�9�9�9:#:c:t:�:�:�:�:�:;C;R;�;�;�;�;<!<A<a<�<�<�<�<�<==+=E=[=n=�=�=�=>$>>>T>n>~>�>�>�>�>??5?Q?a?q?�?�?�?�?�?�?�?�? @    00!030C0W0�0�0�0#131G1w1�1�1�1�1J2�2�2�2�23"3Q3p3�3�3�3�3!4@4[4r4�4�4�455!515A5Q5q5�5�5�5�56Q6r6�6�6�6�6�6A7d7�7�7�7�718X8z8�8�8�8�89:9�9�9�9�9:2:�:�:�:�:�:�:;!;1;A;Q;a;q;�;�;�;�;�;�; <<2<q<�<�<�<�<�<�<=-=@=W=r=�=�=�=�=>!>a>q>�>�>�>�>�>�>�>??!?1?Q?q?�?�?�?�?�?   P  d  00!010A0Q0a0q0�0�0�0�0�011!111A1Q1a1q1�1�1�1�1�1�1�1�122!212A2Q2a2�2�2�2�2�233!313A3Q3a3q3�3�3�3�3�3�344!414A4Q4a4q4�4�4�4�4�4�4"595W5r5�5�5�5�5�566$6>6S6m6�6�6�6�6�67&7@7S7j7�7�7�7848F8t8�8�8�8�8	9$9c9t9�9�9�9�9�9	:A:Q:a:s:�:�:�:�:�:!;1;e;�;�;�;�;�;<<!<A<a<�<�<�<�<=Q=l=�=�=�=>1>Q>q>�>�>�>�>�>�>�>�>??!?1?A?Q?a?q?�?�?�?�?�?�?   `  �   0010Q0q0�0�0�0�01*1<1a1q1�1�13333"3)30373>3E3L3S3Z3a3h3o3v344M4j4}4G5!616a6�6�6�67%7Q7q7�7�7�7�7�78A8a8�8�8�8�8�8�899E9u9�9�9�9:#:3:E:b:{:�:�:�:;%;U;�;�;�;�;<A<a<�<�<�<�<=!=A=c=s=�=�=�=!>1>U>�>�>�>�>o?�?�?�? p  t   A0Q0a0�0�0�0S1a192c2p2�2�2�2Q3�3�3$4U5�5�5�5�5�5�7�78,8G8r8M9f9�:;n;s;�;�; <q<�<=�=�=�=�=>�>??1?I?�?�? �  �   010Q0q0�0�0�01!1A1a1�1�1�1�1�12(2U2u2�2�2�2�23&3:3`3t3�3�3�3�3�3494M4a44�4�4�45E5u5�5�56a6�6�6�6!7A7a7�7�7�7858e8�8�8�89989�9�9�9�9%:Q:u:�:�:;#;=;N;�;5<a<�<�<�<�<�<�<q=�=�=�>�>?=?S?c?�?�?�?   �  �   A0a0�0�0�01E1u1�1�12c2t2�2�2�2�23!3S3j3�3�3	44;4i4�4�4�4�4%5C5f5�5�5j6r6z6�67y7�7�7@8[8�8/9J9R9p9�9�9�9�9C:S:u:�:�:�:�:^;�;�;�;8<�<�<=5=b=�=�=�=8>o>�>�>�>#?3?G?�?�?   �  �   0A0�0:1�1�12
2%2�2�243H3�3�3�3#4<4s4�4�4P5g5�56T6x6�6�67 7n77�7898U8�8�8�8�89C9S9�9�9#:C:�;�;�;<x<S=c=�=�=�=	><>R>�>?=?m?�?�?�? �  �   !0a0�0�0�0/11�1/22�23o3�34_4�4�4O5�5�5=66�67a7�78H8�8�8?9�9�9�98:m:�:�:;[;};�;�;<3<D<n<�<+=n=�=�=�=>>U>�>�>�>)?Y?�?�? �  �   0A0m0�0�0�0!1Q1�1�1�1!2Q2s2�2�2�213]3�3�3�3�3�4�4�45#555T5�5�5�5�5636C6e6�6�677C7]7�7�7�7�7 8888A8r8�89!9W9�9D:�:; ;$;(;,;0;4;8;<;^;Q<�<�<�<�<�<�<�<�<�<�=�=�=�=�=�=>Y>�>�>�>�>�>�>?9?q?�? �  �   �0161s1�1�1C2S2�2�2�23Q3u3�3�3�3�3�34(484s4�4�4�4�45'5:5E5^5w5�5�5�5�56Q6a6q6�6�6�67,7F7j7�7�7�78L8p8�8�8�89Q9i9�9�9�9:4:F:Y:�:�:�:�:
;;-;�;�;�;�;<L<i<�<�<�<�<==v=�=�=:>p>�>A?F?b?~?�?�?�?�?�? �  �   000S0c0�0�0�011�1�1�1#242H2Z2�2�2�2�2�2	3C3T3v3�3�3 4464�4�45t5�56H6�6k7�7T8h89)9e9�9�9:6:;!;;;U;j;�;�;�;<!<�=�=�=�=>C>R>p>�>�>�>Q?�?�?�?�? �  �   0!0A0a0�0�0�0�0181|1�1�1�12%2S2d2x2�2�2�23�3�3�3�344E4^4�4�4�4�4585K5o5�5�5�566E6q6�6�6�6�6717Q7q7�7�7818a8�8�8�8919Q9q9�9�9�9�9:A:x:�:�:�:�:;1;Q;q;�;�;�;<=<Q<f<�<�<t=�=>3>L>r>�>�>�>?>?d?�?�?�?     �   !0A0a0�0�0�0�01!1A1e1�1�1�1�12.2Q2u2�2�2�23!313D3a3�3�3�3!4�4�4�4�45/5k5�5�5686d6�6�6�6�6727J7(838~8�8�8�8�8B9Y;1>J>�>�>�>�>?S?l?  P   1111+1Q1a1{1�1�1�122E2J2a2�2�2�213A3T3�3�3P4�4�4�4�4%5q5�5�5�5x6}6�:   8   ;1�3�4�4�5`6<8@8D8H8L8�8�8�8�8�9�9$:�:;�;<�=�> 0 �   A0�0�0�0151�1�1�1�1�1�1�1�1�2�5
666'6A6�6�6�7868u8�8�89R9v9�9�9�9#:L:�:�:�:;B;q;�;�;<C<S<g<�<�<"=A=b=�=�=>A>i>s>�>�>�>�>?E?x?�?�?�? @ �   (0q0�0�0+1k1�1�122b2�2�23R3�3�34B4�4�4525b5�5�56b6�6�6�6�657�7�78b8�8�8"9b9�9�9B:�:�:�:�:�:6;P;`;�;�;�;<<�<�<=%=1=N=q=�=�=�=>R>^>d>�>�>�>�>?,?0?4?8?<?@?[?d?q?�?�?�?�? P D  010Q0q0�0�0�0�0�0111A1a1�1�1�1�12!2E2a2�2�2�2�2353Q3u3�3�3�344!434A4[4v4�4�4�4�4�455!555a5s5�5�5�5�5�5�56A6Q6c6t6�6�6�6�67$7>7V7p7�7�7�7�7�788!818A8Q8a8q8�8�8�8�8�8�8�8�89/9q9�9�9�9�9�9�9�9A:Q:a:�:�:;;!;1;A;Q;a;q;�;�;�;�;�;�;�;<<4<D<�<�<�<�<�<�<1=A=T=�=�=�=�=>>!>1>A>Q>c>r>�>�>??!?7?_?t?y?�?�?�? `   40e0�0�0�0151a1q1�1�1�122c2s2�2�23Q3a3q3�3�3�3�3�34C4S4u4�4�455$5J5l5�5�5�56"6Y6�6�6�6�6#747N7b7�7�7�7�78c8s8�8�8�89S9c9u9�9�9�9A:Q:a:|:�:�:�:�:�:�:;;!;1;A;Q;a;q;�;�;�;<!<1<A<Q<a<q<�<�<�<�<�<�<�<�<=='=?=O=y=�=�=[>�>�>�>�>�>?L?T?�?�?�?�?�?�? p �   0:0M0R0g0�0�0�0�0d1j1v11�1�1�1�1�12J2X2�2�2�2�2�2�2	3q3�3�3�3�3414A4Q4a4�4�4�4�45'5W5q5�5�5�5�5�56"6@6�6�6�67!7E7a7�7�7�7�7818Q8q8�8�8�8�8�8�8�8�89!919A9a9�9�9�9�9::0:�:�:);D;�;�;<C<T<�<=S=d=�=>c>s>�>?C?S?g?�? � �   #040�0�0#131�1�1�1y2�2�2�2[3�3�3&4A4_4}4�4�4�4g5�5�566Q6o6�6�6�6�6w7�7�738D8�8�8�89c9s9�9:C:T:�:�:;-;s;�;�;<S<d<�<=C=S=�=>>�>�>�>�>3?C?W?�?   � �   0$0�0�011�1�1�1Y2t2�2�2>3�3�3�34!4A4e4�4�4�4555T5r5�5�5�5�56!6�6�6�6�67!7A7Q7q7�7�7�78E8q8�8�8�8�8�8�8�8�89 9%9*9/9G9q9�9�9�9�9�9�9:-:Q:�:�:�:�:�:-;^;�;�;<M<~<�<=!=1=A=�=�=>!>A>a>�>�>�>�>�>?1?Q?q?�?�?�?�?   � �   010Q0q0�0�0�0�0111Q1q1�1�1�12Q2�2�2�2313Q3q3�3�3�3�3414Q4t4�4�4515Q5q5�5�5�5�5616Q6u6�6�6�67!7A7a7�7�738�8�8�8�9�9�9�9C:H:e:j:N;S;�;�;V<[<�<�<N=S=�=�=�=�=   � ,   50`0�566666�8�8�8<�>�>?R?�?�? � �   0R0�0�0�021r1�1�12B2r2�2�2323b3�3�3"4b4�4�4"5b5�5�5B6�6�67R7�7�8�8959e9�9�9�9:1:W:�:3;D;�;!<A<Z<q<�<�<�<�<=!=A=e=�=�=%>U>�>�>�>�>�>�?�?�? � P  80B0G0L0b0n0�0�0�0�0�0�0 11 1,151?1E1M1}1�1�1�1�1�1�1�1�12
22#2/2>2F2]2c2�2�2�2�2=3o3�3�3�3�3�3�3�344414F4Q4g4�4�4�4�4�4�4�4�4�4�4�45E5K5Q5W5]5c5j5q5x55�5�5�5�5�5�5�5�5�5�5�5�5�5 666'6�6�6�6 7f7k7}7�7�7�7X8{8�8�8�8�8�8�8�8�899.94999Q9n9�9�9�9�9�9�9�9�9�9�9�9:::Q:X:{:�:�:;$;+;N;�;�;2<�<�<8=�=�=�=>0>S>v>�>�>J?�?�? � �   0)0L0o0�01C1n1�12�2�23n3�3�3484B4L4o4�4�4�45I5t5�5�5�56;6f6�6�6�67=7`7�7�7�7�78B8e8�8�89S9v9�9�9�92:U:�:�:�:3;s;�;�;<[<�<�<�<"=^=�=�=�=6>r>�>�>*?f?�?�?   � `   	0M0x0�0�01W1�1�1�152`2�2�2�2373b3�3�3�3494d4�4�4�45;5f5�5�5�56=6h6�6�6�6�6�6�677   �  �0�0�0014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�2�2�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�7�7�7�9�9�9�9�9;;;;T;X;l;p;t;|;�;�;�;�;�;�;�;�;�;�;<<<(<,<0<4<8<@<X<h<l<|<�<�<�<�<�<�<�<�<�<�<�< ===$=(=0=H=X=\=l=p=t=|=�=�=�=�=�=�=�=�=�=�=�=>>>,><>@>P>T>\>t>�>�>�>�>�>�>    �  1181@1H1P1\1|1�1�1�1�1�1�1�1�1�12222$2,242<2D2L2T2\2d2p2�2�2�2 3$3H3l3�3�3�3�3�3�3�3�3�3�3�3�3�3�34 4,4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45555$5,545<5D5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5�5�5�5606T6x6�6�6�67,7P7t7�7�7�78(8L8p8�8�8�8 9 9(90989@9H9P9\9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :$:H:l:�:�:�:�:;$;,;4;<;D;L;T;\;d;l;t;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<$<,<4<<<D<L<T<\<d<l<t<|<�<�<�<�<�<�<�<�<�<�<�<�< =D=h=�=�=�=�=>@>d>�>�>�>�>?<?`?�?�?�?�?     �  080\0�0�0�0�0141X1x1�1�1�1�1�1�1�1�1�1�1�122$2D2P2p2|2�2�2�2�2�2�2�2�2�23(3L3l3x3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�45@5d5�5�5�5�56<6`6�6�6�6�6787\7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888$8,848<8D8L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999$9,949<9D9L9T9\9d9l9t9�9�9�9�9:4:X:|:�:�:�:;0;T;x;�;�;�;<,<P<t<�<�<�<=(=L=p=�=�=�=�=�= >(>,>H>h>�>�>�>�> @      0000L0l0�0�0�0�0�01 1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                