MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �V�Z�7�	�7�	�7�	�OX	�7�	�7�	�7�	{yS	�7�	�AU	�7�	�Aa	�7�	�A`	�7�	�AP	�7�	�AV	�7�	Rich�7�	                PE  L ���P        � !
  �       Z�                             �	         @                    0	 ^   �	 (                            �	 �%  `�                                            ̑	 �                          .textbss�                        �  �.text   ��  �  �                   `.rdata  ~�   �  �   �             @  @.data   �D   @	     j             @  �.idata  �
   �	     �             @  �.reloc  �,   �	  .   �             @  B                                                                                                                                                                                                                                                                                                                �������� �/ �� �'W �B� �{� �9� �C� �>� ��� �dg �B. �v � 鰿 �[ ��� �q| �y �7@ �� �S �� �C� �>y �ɩ ��� �/" �� � �pn �Z �6� 鱑 �mc ��. ��z �=� �� �R �� 鉆  鍸 �r �x �� �� �a �6� �r �\l 闉 ��� �m�  騲  �P � �9j  �e 鋯 ��� �U: �� 鋰 �E �q ��  �w�  �Ba �� ���  �c" ��+ �[ �� ��  隚  �� �@m �P" �v� �ak �� �W� �� �]� ��" ��g ���  �I�  �d� ��� ��? �U� �P �7 �E ��> ��+ ��� �r� �BN 鸔 ��/ �>� �YM �O �� �
 �ŉ �@w  �K{  �F0 �� ��� ��  ���  ��1 �H� �N �N� �N� �: �� �� �� �n �k � 遐  �  �7{  �m` �M� �X� �� �N�  ��x �2 �� �: ��) �� �[L �n �`H ��a �y  ��� ��� ��� ��� �^�  �i� �� ��A ��� �E� �Y �{
 �F< �Aa �_ �� �� �]�  ��� 鳿  �z  ��� ��Z �?�  �j  �* �0�  � ��^ ��{  � �g~  鑜 �/ �%n �C� �~� �= �� �� �� 酚  �t\ �� 閔 �A( ��m �W�  ��� �=d �h�  �F �n�  鉻 ���  � �U ���  鐕  �{% �v�  �y �,� ��� ��� �M� �1 �l �� �i� ���  ��� ��l 酡 �D �A ��� �� �& �w�  麫 �} � �� �~� �ټ ��� ��
 �*�  ���  �Ƨ �[�  �fw  �]l �b �0l �B^ ��� �_ ��J �^q �c� �� ��� 骵 �ǫ �`� ��� �Ƹ �a�  �� �7� 馬 � ��� �N ��) � �$� �O� �p� ��� �� �;�  �e  � c �K �g� �'- �B �8�  �s �w �Yp �t+ �/�  �p� � �� �� ��� �l �<�  ��_ �/ � �x�  �e  锳 �O� �� �� ��� �ݪ �k �s �f� ��Q �; 馥 ��[ � �h  �� ���  �� �T- �ό ��  ��  �@� �~ �� �Q�  �[ ��� ��7 �#� ��� �� ��N � ��� �_ �
�  � �P\ �+E �&� �A  �� �7� �7 �� 鈚  �kG ��> �ɖ �Ԫ �1l ��	 ��� ��� �o ��D �Q� �C 駱 邓  ��- ��j �{k �@ �Yj 餔 �_E �� 酠 �0 � �v� ��6 ��� �u ��L �� �" �C �^� �� �b� �� �j� 酑  �� �® ��p � ��  錒 �2  �� 鮗 �t� �Ϊ �	�  養  �� �� �Y �0+ ��w �� �Ak ��@ �w� �� �)� �o# ��Q �D� �&� �:� 鿃  �j �u� �P_ ���  �Ƌ  �}� �l� �m �RP ��  �� ��  ���  �0j � 鏞  � R �' �� �ۂ �6�  �P �M �e� �� �=�  ���  ��  �n� � �$l �J �u �} �0� ��R �V�  ���  風 �_ �k �- �X� �� �&� �i� ��  ��h 鲂 �ը �0� 離 �V� 関 �<� ��  �D� ��L 騇  �Sg �^�  �E_ �Z� ���  �?� �G� ��� �
 ��u �a �L�  �TC �� �g �ρ �ê 龜 �	A �4Z � � �  � �٧ ��� �!� �� �W� �R� ��� ��]  �� �NC �+ �� ��q  �:� �5�  �f� �+u ��X �1( �p  �-� �b� ��  ��� ��� �| �) �T�  �� �j� ��  �`]  �ۅ  ��� ��| �� �'z �b ���  �H �#� �D �M ��� �@ � �er  �@� �E �� �1, �L
 �� �� �!q �g �Cg �� �2� 鄼 �P� ��� �%� ��� ��E �F ��r �lL ��� ��  �[� 鍫 �z� �> �� �) ��� �z�  �E�  �@� ��  �� �q> �, �=� �b� ��  �X�  �3�  �Np �/� � �� �� ��  �@�  ��� �� �!� 鬟 �'7 �2�  �-a  �Ȥ �#F �N� �iJ �� �oG �* �E� �q ���  �s� �� �L@ 鹥 �4� �}�  鲭 �� �;� �	� ��� ���  �:� ��� �pH ��� �� ��3 ���  霭 �� ��  �0� �M� ��� ��� �t  ��  鮿 ��p �@� �: �V �A�  ��L �Ѽ �g ���  �Y ��G ��p �yj ���  �� �0 �� �= �ۋ  �6� �1a �� �[ ��E �� 鸁 �#� ��g  �>� �T�  �O �%� �N ��B ��; �F�  ��� �,� � �h� �]� 鈺 �$� ��< �)�  �� �Y �!l �u�  阔 ��� �ȋ �u �� �#� �: �P 鈼 �s �^N �I�  �Y �Z �Z 鹢 �P ��( �f �: ��� �ǖ  �j �- � � �s� �N� �� �d�  �U� ��� �V � � �k� �F� ��  �,�  �5x �w �� �=5 �� ��� �I� �$� ��N �? �� �з �k  � $ �!� �. �G � �C ��  郘  �H� �� �T �	� �J� �uz ��� �d �V` �}  ��p  �g�  �Q ��� �X� �c> �~�  � �� �/� �jN �U�  鐁 �( �S ��  ��� �A� �r ��Z �f ��5 �n� ��\ �� �
 �J8 ��u �0� ��x �� 锍 ��� �	 �b� ��� �X� � 邡 ��O �D � �*4 �%X �� 饅 �f� �� 鼒 �' �rE �� ��! �� �N� �X� �4W ��  �� �%� � �� �Sa �a  �|� ���  �B �}� ��j  �c� �} �I�  �$�  �: �T �� 頚 �U� �֪ �Q�  �� �L �"
 �M� � 郤 �n' �Ys  �i �� �y �k ��  �[�  �F� ��= �� �W5 �2~  �8� �n �C�  ��� ��� �� �?a �z �EZ �^ �{6 ��� �1% �|I �wm  颳 �� � �� �^�  �Z  �U � �
� �u� � 5 �� ��� �ax ��  �� �( �C� �f ��� �p �	\  �N� �z �ʻ �� �� 馏 閳  �\ ��  駞  �� �� ��� �c� �j  ��: �- ��Z  �� �� �9 �+� �F�  �b �\H �7 �D 齚 ��M �cK � �Y� �c ���  �* �V �" � �&�  �Q�  �� �I ��A �� �(5 �S ��  �p � �� �` �V� �pC �+� �x� �t �|� 駮  �  �- �� �C� �^� �	 �ą �� �
� ��  �@�  �V@ ��� �} �<a  �O �� ��% �О �K �� �^I �� 鿇 ��� �e �p�  �H �Vx �� �f 駐  ��n  �` �h� �� �ԝ � �ĸ �! �Z� �� �`�  �X  �V� ��� 震 ���  �� � � � �f �h �)� �o  �~� 骾 � � � �[ 鼢 ��t �� �7	 ��  �� 騣 ��  �H� �� 鴭 � 麛 �c 逮  �� ��O �y �� �L � �� �hz ��% �[ �� �]W �Ͻ �*n ��9 �� ���  �6[ ��  �ڵ ��� �V� ��� 鸺 �S\ �� �ʥ �� �^ �DK �Uj 鹙 �� �ƞ �1 �l} �f� �@ �2b �X�  ��� 鳴 �iw �$� ��b ���  ���  �C � ��� �g �LN 鷔 �� �Y �X� �Sl �� �i �� �P� 麹 �; �0�  �;� �v� �Q�  鼫  駷 �rw �md 騛  �3- ��@ �j �N� �& ��� �� �g �[j 鶸 �v �	� �q �[ �M� �H� �J �? �[� �Ax � �*r ��9 �� �k �f� �!` �� �� ��_ 靳  �( �Cs ��  �� ��y �y� �x� ��  �a ��� 鶴 �T� ��N 駙 �� �]� �8	 �~  �� �%{ �$ �h  ��� ��� �� ��q ���  �a�  鬫 ��h �"�  ��� �X+ ��= �NM �Y� �]G 鿷 �
7 �� �� �{� �&  �m ��w 釄 ��s �w� ���  郆  �>q �	d �d� ��  �# �^ �8 �= �� �a �M �� �bT �L �j  ��I �hG �	� �D� �O�  ���  �c ��� 鋒 �ֶ  遶  �ܥ  �', ��r  �� � ��  �n �_� �? �� �� �� �PX � �� �A� ��B �g �2� �mQ  �[ ��� ��: ��C �D� �G� �A �� �= ��+ �� ��B �G �� �� �/� �(f ��N �~�  �	 �B ��l  �J� ��� � �  ��  ���  ��  ��� ��C �"�  锔 �� �3| � �� �� 饍 �PD ��w �pS �# ���  ���  �q 野 �2Q �s ��|  鳸 �Y �y� ���  鿘  �đ �j� ��. ��0 �� �4� ��  ��� �B� ��{ �V �� �>� �	�  �4: �Ϡ �zi �jc �G �00 �& �  �� ��  �b�  ��  � � �Q� �I� ��s �t� �Op �J �E�  �Ц �[�  ��- �� �e ��\ �b� �a � ��  �>�  �i�  餼 ��  ��k �� ��= �= 馺  �q9 �y� �- ��D �-� �� �< �>�  �y � �_� �? �� �� �;� �� �ݕ ��� �gK �"� �) ��Y �c�  �Ζ ��A �t�  �� �
L �E� ��e ��0 �ց  �ѯ  �w �O� �� 靏 �� �� �n� �  餅 ��> �� �o ��  �y� �V� �aI �� �'�  �� �my �= �� �� ��l �� ��� �z� ��  �� �> 鶿 �� �,� ��5 �m �� �HQ �N� ��  �� �t� ��� �z� �a  �� �yU ��x �u  �`  �3 �B� ��� ��� �$ �� �G� ��� 鑕 �z� �%� ��� 鋆  �jm �u �<B �g� �Ҍ �mP  �� �I � ��  �T� ��� �l �� ��0 � � 閜 ��� �� 释  �r� �͎ � 韔 �R� �B �D�  �?u  � �& ��  �`  邯 ��) �`� �7_ � 驏 � ��� ��� �{ �$: �� ��> ��' ��� 髣 ��  �q� �� �] �R] �͘ �� �s� ��v ��$ ��  �;� �*� �E�  ���  ��� � ��Y � �w�  �|� ��  騉  �c�  �N� �Ib �< �� ��\ �<] �p�  �AU �� �n �\� ��u �< �}7 ��� 飆 ��  �[  �j �� � ���  ���  �� 醔  �az  �� �� �B� ��i �X�  ��
 �~�  �t� �4` ��� ��� 鵼 鐵 �[�  ��y  �� � � �'�  �r�  �OO �^� �s ��j �= �� �$ ��k 鵝 �' �{! ��� �!� �,� 鷈  ��  �g� �� �ҷ �3S �L� �tb  ��I �
� �T � � � �1> �� ��  �< �,s �� �s# �^ �� �y8 ��� �� �Ղ ��t  �l ��S �Ѡ �\d �K� 釸 �L �hn �c& �$ �� �d� �� �: �L ���  �-6 �V �+� �,. �, �b� �H6 �H� �X �.}  �9u  �� �O� �� �fF �3I ��l 閷  ��  ��c  ��  �8� �_ �� ��  �#0 ���  � �� �  �U]  ��k �g �\ �Y �) ��  ��  �=� �h 雮 �3 � 鄔 �o ��� �ȷ � � �{� �H  �
 �� �1x ��� ��� �1 �s� �8 �s �L �/{  �:r  �
H �� ��X �&�  �!�  �<| �7�  �"� �� �c �}  �F  �� 餕 �� �Zq �k: � | �r �&� ��� �<H �] �X �MD �.T �S �N
 �	�  �d# �?� �ڜ ��  �0� 黺 �c� �� �? 鴥 �r� � �Ȩ  �� �[ �y�  �� �S �� 鯎 �� ��  鶙 �KO �L�  �� �rx  � �� ��� �� �	 �T �� �~  �O �� �o �] � �\� 飏 �_� �� �H �ê �n�  �\ �4�  �^  �Z0 ��� �К �+�  �^d ��k �� �B �� �6 鸋 ��f �N�  陼  �4� �o� ��� �: �@� �� �V �- � �ˆ �r| �}� �x� �S� 鮓 �]: �$ 鏭 �
$ ��  ��W �� �� �� �� � ���  �M] 鈖 郴  �΃ �� 鴑  ��}  �(g �EK �� ��= �ʍ �T �<X �G� ��z �3 �� �CT �	 �i�  ��@ ��p ��! �< ��6 ��� �&� ��x �|� �'� �r�  �]�  �[f ��� �@ �� 鲌 �J ��
 �r1 �P� �� �� �Y �,� �G�  �2� ��  ��F  铐 �^�  ��X  �U  �Ì ��k �e� ��� �D �� �1� �\s  �"� �V� �� �) ��z  �� �| �\ �� �N �{. �T �� �v� �� �l~ �G�  �: �`~ �e �) � �	h �H  鍋 ��r �d ��S �+�  �X 铋 �<�  �W{  锘 �� �xx �� �~K �W� 雳 �� �u �E� �P�  颓 �3" ��� �� �ǝ  �a� �L �Ȯ �Q �� �٥  �� �) �v �d �@� �K�  �� �l  ���  �� 鷔 �� �� ��6 �^� �)�  �?� �� ��: �%{  預 �{v �� �1� �?3 ��  ��1 �~ ��� �3� ��� �ɴ  ��? �� �� 鍀 逝 ��D �A �/ �|~  駤 ��  ��� �� ��i  �� �iI  �K� �O# �z� � � �  ��� ��; �! ��: ��  �t� ��A �K �K �nT �� �D ��3 �ha �z  �p| �K� � �A@ �|�  �: �ka �Mx  �U  �5� 鎛  �If  �T\  �Z ��Q �5| �P�  鵉 ��� �4 �ܞ ��� ���  �b �h: �L �� ��A ��% �@5 �
� ��� �`P ��6 ��3 �і  鼉 ��  �K  �܁ �H� �� �>{  �E� �(� ��0 �)� �X# �0Y � �f	 �� �lk  �F3 �B� ���  ��� �V9 �~ �� �D� ��  隆 �� �G �[� ��q �a� �� �g� �B� �ݿ �h�  �sq  � �q� �H� ��� �*� �� �@ ��% � �� ��# � �b�  �g �8�  飘 ��  鹪  �d� ��  �e ���  �p�  ��K �כ �#� �,�  �g� �?  鍁 �ع �� �& �ɬ �. �?< �z�  ��c  �  �[6 ��� ��@ �ܯ  ��� �R� �}U  �XJ  �/O �Ϋ �Yy �X �� ��� �� �p �E � � �_� ��` ��) ���  �H�  �� �8 �. �J �  ��  �K  � �;�  �!� �e- �\�  ��� ��L �MV �"� �# �, ��  �� �5 �ھ �u�  � � �u� �&8 �q �j �� �� �l �h3 �SQ �~; 陁 ��G �� �"S �g3 �C ���  �vw  鞜 �
 �� �2? �R �}R �c' 龦 鹻 �t�  � ��4 �E� � f 鰁 鈋 �8 �� �YF ��@ �� 鈹 鳓 �5 ��  �` 麪 �M �	� � � �� �?  ��� ��  ��� � �]�  ��w  �0� �b~ �;� �d�  �� ��� �7� � 颎 �~ �� �J� �G9 �b�  �/� ��8 �#�  �Nj  � �dH  ��F ��: �e �P{ ��S �vv  �!J �� �� ��  �� ��a ��  � �{ 餠  �� �z� �� �� ��  ��  �l 鬃 �w�  �� ��{ �Є � �F ��M �� �ߧ �* �% � t  � �!� 驩 �5 ���  �� �j� �(c �u  �_ ��[ �T�  ��  �� �A� � � �K� ��F �� �L@ �� ��t �=� �� �� �rq �v �dt ���  �b� �� �@�  �K� �� �)� �|' �W� �"� �� 鼃 �� �" �� �T �o�  �V �%�  ��� �� �  ��� �<v �� ��  �=�  ���  �� � � 錿 �q �/� 銵  �' � . �+M  鳵 �� �D ��~ �" �=� �x�  ��� �~I �	$ �o� �o� �m �uG �#� �+O ��  �v �p� �8 ��  �h �� �ɾ �t� �j �% �?� �� ��  �: ��n 鶾 �a � ��* �D �+ �E� �� �� �n �\ �l �+ �Z �> �
� �7n 鑤 �� �g�  ��� �x  �X� 郔  酋 �� �4# � �Jh 雃 �@ ���  �c  �� �|5 ��e  �D� ��6 ��� ��  �.�  �ں �. �u1 �w ��� �P� 鑁 飋 ��  �� ���  �2�  ��  �u �+ � � �T �, �4� �� ��� �KR �I ��� 餼 �W�  閂 �� �hM �c� �~r �)8 � 鿚 �� �u\ � �  �;� �� �qT ��� �W� �2O �]�  �^ �'� ��
 �ə  �� �/+ 骄 � �� �+� ��N �a�  ��  �� �2 �=�  鍮 ��� �Vp � � �?� �
 ��X � � �� �Y ��f  �*@ �� 邩  ��  �� ��  �� ��v �dJ  �'� ���  ��6  �5� �<3 �oY �m� �%M �<� �o  �� ��  �� �� �y� ��f �� �zb �� �� ��x �> �ь �L� ��t ��l ��' ��9 �� 龦 ��X ��D �oA �� �H� �P� �ۿ �6# �7  �v� �I  �� �� ���  �M/ �~�  ��� �d�  �� ��+ �%  �p 雯  ��! �� �Lm �! 钂 �k  �L �c�  ��X �+ �i �? ��� �@ �@m  鐞 �6  �V �) �� �� �� �� �#�  �>] �z �d[ �&r �*� ��  騗 �5 �" ��_ �$ �3 �c �� �x�  �%~ �,� �y�  �4� ��1 �� ��0 ��f �W �6p  �Q�  �<�  駅 �B� �m- �� �3 �.�  �#� ��t  �� �
� �� �`` ��B �&�  � �<� �G �Rl ��N  � ��� �^ �Ie �� ��� ��}  �~ ��  ��1 ��b  ��� ��} �O� ��� �] �� �C�  �A: � �� �f �Z ��� ��5  �F> � ��# �� �z� �� �]  �h� ���  �n� �٤ 鄮  �W �t} 鵑 �p �˴ �W �Q �Lp �w�  �� �[ �(�  ��; �� 鳵 �� �f �J@  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@SVW�E���Ex�M�U�EE�E��_^[��]� ������������������U���@SVW耰���   _^[��]�������U���DSVW�E�E��}�t��@Z	������   _^[��]������������������U���@SVW_^[��]�����������������U���LSVW�E�    ��M������E�} t^�EP�MQ�M负���M������E��} t2�}� t,j �EP�MQ�UR�E�P袡�����E�} t	�E�E�E��E����E�둋E�_^[��]��������������������������������������U���DSVW�M��TZ	���   �M��B(��_^[��]�����������U���DSVW�M��TZ	���   �M��B4��_^[��]�����������U���HSVW�E�    ��M������E�} t*�EP�M������E��E�;Eu�E����E��} t��ŋE�_^[��]��������������������������U���pSVWj h���M������E�P�M��`����M��ٛ���E�    �E�    j h���M������j �M�� ���P�E�Ph��j j �Ι����PhD� �N������E��M�胛���M��4����E�_^[��]���������������������������������������������U���DSVW�M��E�P�TZ	�Q�B�Ѓ��EPj��MQ�U�R�TZ	�H�Q�҃��E�_^[��]� ���������������������U���DSVW�M��E�P�TZ	�Q�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�� _^[��]���������U���HSVWhЮjEhH_	j�E������E��}� t�M������E���E�    �E�_^[��]���������������������������U���DSVW�M��M�訞���E�� D��E�_^[��]����������U���dSVW�M��EP�M�������E��}� u�E��k�M� ����E�jh�  �M��N��������$�����$�����$�M�蘧��Ph�  �M������E��x t�E���P�K������E�_^[��]� ��������������������������������������U���DSVW�M��E��E��E��E�X�E��E�X�E�_^[��]� ��������������U���DSVW�M��EP�MQ�TZ	�B�M��P4��_^[��]� ������������������U���DSVW�M��EP�MQ�TZ	�B�M��PH��_^[��]� ������������������U���DSVW�M��E�P�TZ	�Q@�B,�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M��T����E��x t�E���P������_^[��]� �����������������������U���LSVW�M��EP�MQ�UR�M������E��}� u�E��U�E�P�M������u3��A�E��x t�E��H裫���耚���M��A�}� t�E��HQ�M������u3���E�_^[��]� ������������������������������������U���HSVW�M��EP�MQ�M��*����E��}� u�E��I�E�3Ƀx ��Q�M�֓����u3��,�E��x t jj h�� �E��HQ�M�v�����u3���E�_^[��]� ������������������������������������U���PSVW�M��EP�MQ�UR�M��ӗ���E��}� u�E��V�E�E�E�E��}�t�}�t�}��F t"�0�EP�M�Q�M�������E�P�M�������EP�M�Q�M�輝���E�_^[��]� �����������������������������������U���   SVW�M��M肾����P�M觰��� �E��E������E���D�����D������  ��D�����D�����  ��D����$�2j jjj?�M����P�������E��E��  ��  �E�    j jjj?�M�ĩ��P躙�����E��  �  j jjj?�M藢��P蕙�����E��E��  �t  �E�    j jjj?�M�h���P�f������E��  �H  �M�菸��j��H���P袵����P�M��:�����H����������d����u���Pj�Ȓ����Pj j�M��A����EЍ�d����{����}� ��   �E��x u�[����M��A��E��H�d����E��x uj�o�����P迱�����j j��E�P�M��I�Ǒ���Ẽ}�tj�Ĭ�����E���P�������H�����E�j jj@j@�M�諔��jjh   �E�P�M��I観���E���P蠔�����E��MȉH�M��������E��x t�E���P�u������}� |6�M�ܙ���EċE�P��t���Q�޶����P�U�R�M�������t����U���_^[��]� �I (0P0�1�/�/�1�1|0�1��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���DSVW�M��E�P�TZ	�Q�B�Ѓ��E�_^[��]����������������������U���PSVW�EP�M�Q�TZ	�B�H(�у�P�M輷���M������E_^[��]��������������������U���DSVW�M��E�P�TZ	�Q�B�Ѓ��E�P�MQ�TZ	�B�H�у��E�_^[��]� ��������������������������U���DSVW�M��EP�MQ�TZ	�B�M��P8��_^[��]� ������������������U���DSVW�M��TZ	���   �M��B4��_^[��]�����������U���hSVW�M��M�Z����E�j jj?�M�r���P�ʫ����P�E�P�K�����Ph�  �M�������M��Đ��j jj?�M�0���P萫����P�E�P������Ph�  �M�达���M�芐��_^[��]� ��������������������������������������������U���   SVW�M��E��M��E��x tU�E��8 t�E���M�E�P�M��I������E��H�>����E��E�    �E�    �M��o����E�M�萷���E��m�E���M�}� u�Œ���E�j jj@j@�M�肐���E�PhD� �n�������t�E�P�M��	菜���E��H�M��E��H�M�E��H�M�E��H�M�}� �  �M躕���E�j h�  �M�茧���E܃}� �  ��D���踭��Ph�  �E�P�M���������M��:����E����M��)����E����M������E��M��	����E��E虃�����E܉E�jjj?�M�?���P蟩��������   �E�    �	�E����E��E�;E�}k�E��E��E�   �	�E����E��E�;E�I�E�E�+E��E��E�P�M�Q�U�R�E�P�M�Q�M������}� th�   �E�P�M�Q�U�R�M�������jjj?�M裢��P�����������   �E�    �	�E����E��E�;E�}k�E��E��E�   �	�E����E��E�;E�I�E�E�+E��E��E�P�M�Q�U�R�E�P�M�Q�M��`����}� th�   �E�P�M�Q�U�R�M��I�����3������E��M��H�E��M�H�E��M�H�E��M�H�E��M��E�@   �
�E�@    _^[��]� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���DSVW�M��E�����E����X�E����X�E�_^[��]��������������������U���DSVW�M��EP�MQ�TZ	�B�M����   ��_^[��]� ���������������U���\SVW�M��EP�MQ�U�R�TZ	�P�M����   �ЋM���P�Q�P�Q�P�Q�P�Q�@�A�E_^[��]� ������������������������������������U���DSVW�M��E�P�TZ	�Q�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�Q�B�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�H��  �҃�_^[��]� ����������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�B��  �у�_^[��]� �������������������U���LSVW�M��EP�MQ�UR�EP�MQ�M�货���E��}� u�E��2�E�E�E�x t�E��P�Պ�����E��H�����M�A�E�_^[��]� �������������������������������U���DSVW�M��M������E��t�E�P�z������E�_^[��]� ����������������������������U���DSVW�M��M��Χ���E�� <��E�_^[��]����������U���DSVW�M��M��y���_^[��]����������������������U���DSVW�M��M��2���_^[��]����������������������U���DSVW�M��M������E��t�E�P蚏�����E�_^[��]� ����������������������������U���DSVW�M��M��ŉ���E�� ��E�_^[��]����������U���DSVW�M��M�裔��_^[��]����������������������U���DSVW�M��M��R����E��t�E�P�������E�_^[��]� ����������������������������U���DSVW�} t�E�E���@Z	�����E��M�Q�UR�EP������_^[��]������������������U���DSVW�M��E�� _^[��]���������U���DSVW�M��E��     �E��@    �E��@    �E��@    �E�_^[��]��������������������U���DSVW�M��M�蠒��_^[��]����������������������U���PSVW�M��E��x t�o�E��8 t �E��Q�TZ	�B<�H�у��E��     �E��x t>�E��x t+�E��H�M��U��U��}� tj�M�茗���E���E�    �E��@    _^[��]������������������������������������U���DSVW�M��M��n����E��t�E�P��������E�_^[��]� ����������������������������U���dSVW�M��E�P�&�����P�M��.����E��M������E�_^[��]���������������������������U���LSVW�M��E��x uTh8��|@	��PhH_	j�B������E��}� t�MQ�M��i����E���E�    �U��E��B�E��x u3��H�E��x t�E�3Ƀ8 �����0�EP�TZ	�Q<��Ѓ��M���E��@   �E�3Ƀ8 ����_^[��]� ������������������������������������������������������U���DSVW�M��E��@   �TZ	�H<�Q�ҋM���E�3Ƀ8 ����_^[��]���������������������U���DSVW�M��E��x t�   �+�E��x u3���E��HQ�U��P�TZ	�Q<�B�Ѓ�_^[��]�����������������������������������U���DSVW�M��E��8 u�TZ	�H���EP�M��R�TZ	�H<�Q�҃�_^[��]� �����������������������������U���@SVW�@Z	����_^[��]�������U���@SVW�EP�@Z	�g���_^[��]�������������������U���hSVW�EP�@Z	�7���P�M��Ǩ��j h���M��6���j �E�P�M�Q�M��F���������E��M������U���t�M覤���M��ʂ���E�9j�E�P�M������j�j��EP�M�Q�M������E�P�M�I����M�菂���E_^[��]�������������������������������������������������U���DSVW�M��EP�MQ�UR�TZ	�P�M��B@��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�B�M��PH��_^[��]� ������������������U���DSVW�M��EP�MQ�UR�EP�TZ	�Q�M��BL��_^[��]� ��������������������������U���|SVW�EP�@Z	臮��P�M�����j h���M�膦��j �E�P�M�Q�M�薢��������E��M��2����U���t�M������M������E�   j�E�P�M��F���j�j��EP�M�Q�M��:���j h���M�����j �E�P�M�Q�M��!���������E��M�轀���U���t�M聢���M�襀���E�9j�E�P�M��Ԏ��j�j��EP�M�Q�M��Ț���E�P�M�$����M��j����E_^[��]����������������������������������������������������������������������������U���   SVW�EP�@Z	����P�M�褥��j h����t�������j �E�P��t���Q�M������������s�����t��������s�����t�M�t����M�����E�   j�E�P�M��č��j�j��EP�M�Q�M�踙��j h���M�菤��j �E�P�M�Q�M�蟠��������E��M��;���U���t�M������M��#���E�   j�E�P�M��O���j�j��EP�M�Q�M��C���j h���M�����j �E�P�M�Q�M��*���������E��M���~���U���t�M芠���M��~���E�9j�E�P�M��݌��j�j��EP�M�Q�M��ј���E�P�M�-����M��s~���E_^[��]���������������������������������������������������������������������������������������������������������������������U���   SVW�EP�@Z	�����P�M�脣��j h����`�������j �E�P��`���Q�M�������������_�����`����}����_�����t�M�T����M��x}���E�  j�E�P�M�褋��j�j��EP�M�Q�M�蘗��j h����t����l���j �E�P��t���Q�M��y����������s�����t����}����s�����t�M�О���M���|���E�   j�E�P�M�� ���j�j��EP�M�Q�M�����j h���M�����j �E�P�M�Q�M������������E��M��|���U���t�M�[����M��|���E�   j�E�P�M�諊��j�j��EP�M�Q�M�蟖��j h���M��v���j �E�P�M�Q�M�膝��������E��M��"|���U���t�M�����M��
|���E�9j�E�P�M��9���j�j��EP�M�Q�M��-����E�P�M艡���M���{���E_^[��]�������������������������������������������������������������������������������������������������������������������������������������������������U���@SVW�EP�TZ	�Q<�B�Ѓ�_^[��]������������U���   SVW�E�    j h����l�������P�J~�����E���l�����z���}� u3���   �E�    �E�P�M������E�P�M�Q�M��K�������   �}���   �M������E�}� t:�EP�M��>����M�Pj�M�Q�M�蘝���M����}����tǅh���   �
ǅh���    ��h���������E���t�e���M��z���M���t�e���M���y���������t�E��E���=����E�_^[��]����������������������������������������������������������������������������������������U���DSVW�M��EP�M���x�������_^[��]� ������������������������U���DSVW�M��EP�TZ	�Q�M��Bx��_^[��]� ����������������������U���DSVW�M��E�P�TZ	���   �BT�Ѓ�_^[��]����������������������U���TSVW�M��EP�MQ�U�R�TZ	�P�M����   ��P�M�C����M��x���E_^[��]� ������������������������U���   SVW�E�    �} u6j h����p����j���P�{�����E��p����#x���} u3��   �E�    �EP�M��?����E�P�M�Q�M�襓������   �}���   �M��>����E�}� t:�EP�M�蘙���M�Pj�M�Q�M������M����]z����tǅl���   �
ǅl���    ��l����U��E���t�e���M��ow���M���t�e���M��[w���U���t�E�E��2�+�}�u%�}� t�EP�M��&x������y����t�E�E�������E�_^[��]�������������������������������������������������������������������������������������������U���DSVW�M��E�P�TZ	���   �BH�Ѓ�_^[��]����������������������U���PSVW�} u3��   �EP�M�菀���E�    �E�    �E�P�M�Q�M�������tT�}�t�}�u"�EP�M��~��P�g�������t�   �*�$�}�u�EP�M���v�����x����t�   ��3�_^[��]������������������������������������������������U���@SVW�TZ	�H<�Q��_^[��]��������������������U���DSVW�M��E��@    �E��     �E��@    �E��@   �E�_^[��]��������������������U���DSVW�M��} u�4�} t�EP�M踢��� �} t�EP�M��x����E�P�M�x��_^[��]� �������������������������������U���DSVW�M��EP�TZ	���   �M��B@��_^[��]� �������������������U���DSVW�M��EP�TZ	���   �M��BD��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q@�M��Bd��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q@�M��Bh��_^[��]� ����������������������U���DSVW�M��EP�MQ�TZ	�B@�M��Pl��_^[��]� ������������������U���DSVW�M��EP�MQ�TZ	�B@�M����   ��_^[��]� ���������������U���DSVW�M��EP�TZ	���   �M����   ��_^[��]� ����������������U���DSVW�M��EP�MQ�TZ	���   �M����   ��_^[��]� ����������������������������U���DSVW�M��TZ	�P@�M��Bt��_^[��]��������������U���DSVW�M��TZ	�P@�M��Bx��_^[��]��������������U���DSVW�M��EP�TZ	�Q@�M��B|��_^[��]� ����������������������U���DSVW�M��TZ	�P@�M����   ��_^[��]�����������U���DSVW�M��TZ	���   �M��Bt��_^[��]�����������U���DSVW�M��EP�TZ	�Q@�M����   ��_^[��]� �������������������U���DSVW�M��TZ	�P@�M����   ��_^[��]�����������U���DSVW�M��EP�TZ	�Q@�M����   ��_^[��]� �������������������U���DSVW�M��EP�MQ�UR�EP�TZ	�Q@�M����   ��_^[��]� �����������������������U���DSVW�M��EP�MQ�UR�TZ	�P@�M����   ��_^[��]� ����������������������������U���DSVW�M��EP�MQ�UR�TZ	�P@�M����   ��_^[��]� ����������������������������U���DSVW�M��EP�MQ�TZ	�B@�M����   ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�B@�M����   ��_^[��]� ���������������U���HSVW�M��E�P�TZ	�Q@�B�Ѓ��E��E�#Et�E��#E��E��	�E�E�E��E�P�M�Q�TZ	�B@�H�у�_^[��]� ����������������������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�B@�HL�у�_^[��]� ������������������U���DSVW�M��E�P�TZ	�Q@�BH�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q@�B�Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�M�Q�TZ	�B@�H�у�_^[��]� ������������������U���DSVW�M��EP�MQ�U�R�TZ	�H@�Q�҃�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�B@�H �у�_^[��]� ������������������U���DSVW�M��EP�MQ�TZ	���   �M��P��_^[��]� ���������������U���DSVW�M��EP�MQ�UR�TZ	���   �M��B��_^[��]� ����������������������������U���DSVW�M��EP�MQ�UR�TZ	���   �M��B ��_^[��]� ����������������������������U���DSVW�M��EP�MQ�UR�EP�TZ	���   �M����   ��_^[��]� ��������������������U���DSVW�M��EP�MQ�UR�TZ	���   �M���D  ��_^[��]� �������������������������U���DSVW�M��E P���E�$�MQ�UR�EP�MQ�TZ	���   �M����   ��_^[��]� �����������������������U���DSVW�M��EP�MQ�UR�EP�MQ�TZ	���   �M����   ��_^[��]� ����������������U���DSVW�M��TZ	���   �M��B$��_^[��]�����������U���@SVW�TZ	�H@�Q0��_^[��]��������������������U���@SVWj�EPj �TZ	�Q@�B4�Ѓ�_^[��]������������������������U���@SVWj�EPh   @�TZ	�Q@�B4�Ѓ�_^[��]���������������������U���@SVW�EP�MQj �TZ	�B@�H4�у�_^[��]����������������������U���@SVW�TZ	�H|���_^[��]���������������������U���@SVW�E�8 t�E�Q�TZ	�B|�H�у��E�     _^[��]�������������������������U���@SVW�TZ	�H|�Q ��_^[��]��������������������U���@SVW�E�8 t�E�Q�TZ	�B|�H(�у��E�     _^[��]�������������������������U���@SVW�TZ	�H@�Q0��_^[��]��������������������U���@SVW�E�8 t�E�Q�TZ	�B@�H�у��E�     _^[��]�������������������������U���@SVW�EP�TZ	�Q@���   �Ѓ�_^[��]�������������������������U���@SVW�E�8 t�E�Q�TZ	�B@�H�у��E�     _^[��]�������������������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�BH��d  �у�_^[��]� ���������������U���@SVW�EP�MQ�UR�EP�TZ	�Q �BH�Ѓ�_^[��]����������������U���DSVW�}qF t�1�E�E��}� u�#�EP�M���j���E�P�MQ�M�0m�����֒��_^[��]���������������������U���DSVW�M��EP�MQ�TZ	�B�M��Pp��_^[��]� ������������������U���DSVW�M��TZ	�P@�M��BT��_^[��]��������������U���DSVW�M��EP�TZ	�Q@�M��BX��_^[��]� ����������������������U���DSVW�M��EP�MQ�TZ	�B@�M��P\��_^[��]� ������������������U���DSVW�M��TZ	�P@�M��B`��_^[��]��������������U���@SVW�EP�MQ�TZ	�B��T  �у�_^[��]���������������������U���@SVWh��hE  �M�k���������Ph��hE  �M�yk���������P�TZ	�H��T  �҃�_^[��]��������������������������U���@SVW�E�TZ	�TZ	� _^[��]������������������U���DSVW�M��   _^[��]� ������U���DSVW�M�_^[��]� �����������U���DSVW�M��   _^[��]� ������U���DSVW�M��   _^[��]� ������U���DSVW�M��   _^[��]� ������U���DSVW�M��   _^[��]� ������U���DSVW�M�_^[��]� �����������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�3�_^[��]� ���������U���DSVW�M��   _^[��]� ������U���DSVW�M��   _^[��]� ������U���DSVW�M��   _^[��]� ������U���@SVW�E�M�H4�E�@��E�@8u��E�@<\��E�@@7��E�@Di��E�@H��E�@L4��E�@P���E�@l[��E�@X��E�@\��E�@`d��E�@d3��E�@T.��E�@h���E�@p ��E�@t8��E�M�H �E�M��E�M�H0�E�M�H(�E�@,    _^[��]�����������������������������������������������������������������U����   SVWj h�   ��`���P�������j �EP�MQ�UR�EP��`���Q蓆�����E �E�h�   ��`���P�MQ�URj��u����_^[��]�����������������������������������U���@SVW�EP�M���   Q�UR��e����_^[��]�����������������������U����   SVW�M��c���M���E��8 u��   �EP�� ����Kc��j hб��X���螅��P��<����-c��j j��� ���Q��<���R��h���P�d����P�M�Q�t����P�U�R�t����P�E����]��������؈�����M��Rh���M��Jh����h����?h����<����4h����X�����_���� ����h���������t�E�P�`�����E�_^[��]� �������������������������������������������������������������������������U���DSVW�M��EP�q�����M���E�_^[��]� �����������������������U���DSVW�M��E�P��_����_^[��]�����������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U���  SVW�M��} u0�E��M���P�Q�P�Q�P�Q�P�Q�@�A�E�  �EP�M�Q�U�R�b�����E��HP�������������^  �������$�`nj j �E���@�$�M����$�UR�E���P������Q��z����P�UR�E�P�����Q�Eb����P��(���R�M�������M�P�U�H�M�P�U��H�M�P�U���  �E�P�M���A�$�U����$�EP�M���Q��@���R�Qz����P�EP�M�Q��X���R��a����P��p���P�M�]����M�P�U�H�M�P�U��H�M�P�U��}� ��  �����$�����$�����$�������Oj��P�EP�M�Q������R�Ha����P������P�M�5p��P�MQ�U���R�E�P������Q�W����P������R�	a����P�� ���P�M��o��P�����Q�Nt����P��0���R� t����P�E�P��k�����EP�M�Q��H���R�`����P�E�P�MQ�U�R��`���P�`����P��x���Q�M�o��P������R�W����P������P�M�f��P������Q�s����P������R�s������MȋP�ŰH�MЋP�UԋH�M؋P�U�j j �E���@�$�M����$�U�R�EP�M�Q������R��_����P�����P�M詄����M�P�U�H�M�P�U��H�M�P�U��w  �E�@��������D{8�EP�� ���Q�M�e����U�H�M�P�U�H�M��P�U�@�E��q�E�P��P���Q�M�jl�����@�$�U���B�$�E��� �$��8���� h��P��h���Q�M�@e����U�H�M�P�U�H�M��P�U�@�E��  j �E���@�$�M����$�UR�E���P������Q�?w����P�UR�E���0P������Q�^����P������R�M�jZ����M�P�U�H�M�P�U��H�M�P�U��E���0P�M�Q������R��q����P������P�q����P�M����AH�$������R�b����P�E���0P�����Q��T������U�H�M�P�U�H�M��P�U�@�E��  j�EP�M���0Q��(���R��]����P�M�\r���E��HH�]��E���������Dz	���]��EP�M���0Q��@���R�]����P��X���P�M�l��P�MQ��p���R��p������M�P�U�H�M�P�U��H�M�P�U����]���E��$�E�P�k������$�Nd�����]��E�P������Q�Yp����P���E��$������R�ha������M�P�U�H�M�P�U��H�M�P�U��E��u����$��q���$�݄�������M��]�EP�M���0Q������R�\����P������P�M�k��P�M�Q������R�S����P�� ���P�M�b����M�P�U�H�M�P�U��H�M�P�U��EP�����Q�*j����P�U�R�EP�\�����E_^[��]� �gdh�jxk~l����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@SVW�E�]����Au�E��E_^[��]������������U���@SVW���E�$�)m����_^[��]����������������U���@SVW���]����Az
�8��+��(��]����u������E�$��{����_^[��]����������������������������������U���@SVW�E�M� �I�U�E�B�����$�M�U�A�
�E�M� �I����$�U�E�B�H�M�U�A�J����$�M��a���E_^[��]������������������������������������������U���@SVW�E�M� �	�U�E�B�H���M�U�A�J�����$�4X����_^[��]�����������������������������U���@SVW���E�$�}m ��_^[��]����������������U���HSVW�E�M� �	�U�E�B�H���M�U�A�J�����$�W�����]��E���������Dz�����$�M�%b���E�?���u��]��E�@�M����$�M�A�M����$�U��M����$�M�`���E_^[��]��������������������������������������������������������U���DSVW�M��E��E��E��E�X�E��E�X�E�_^[��]� ��������������U���@SVW�E�@�M���$�M�A�M���$�U��M���$�M��_���E_^[��]��������������������������U���@SVW�E�M�@�A���$�U�E�B�@���$�M�U�����$�M�[_���E_^[��]����������������������������������U���@SVW�E�M�@�a���$�U�E�B�`���$�M�U��"���$�M��^���E_^[��]����������������������������������U���@SVW�E�M�@(�	�U�E�B@�H���M�U�AX�J�����$�E�M�@ �	�U�E�B8�H���M�U�AP�J�����$�E�M�@�	�U�E�B0�H���M�U�AH�J�����$�M�(^���E_^[��]�����������������������������������������������U���@SVW�E�M�@(�	�U�B�E�M�@@�I���U�E�BX�H�����$�M�U�A �
�E�@�M�U�A8�J���E�M�@P�I�����$�U�E�B��M��U�E�B0�H���M�U�AH�J�����$�M�G]���E_^[��]����������������������������������������������U���   SVWj �M��IO���E�M�@8�IX�U�E�BP�H@��M�I�U�E�BP�H(�M�U�A �JX��E�H0���M�U�A �J@�E�M�@8�I(��U�JH���]��E���������Dz�M��m���E�s  ���u��]��E�M�@�IX�U�E�BP�H��M�I0�U�E�B�H8�M�U�A�J@��E�HH���M�U�AP�J@�E�M�@8�IX��U�
���M��]��E�M�@�I(�U�E�B �H��M�IH�U�E�B �HX�M�U�AP�J(��E����M�U�AP�J�E�M�@�IX��U�J���M��]��E�M�@8�I(�U�E�B �H@��M�	�U�E�B@�H�M�U�A8�J��E�H���M�U�A�J �E�M�@�I(��U�J0���M��]��E�M�@8�IX�U�E�BP�H@���M��]��E�M�@P�I(�U�E�B �HX���M��]��E�M�@ �I@�U�E�B8�H(���M��]ȋE�M�@@�IH�U�E�BX�H0���M��]ЋE�M�@X�I�U�E�B(�HH���M��]؋E�M�@(�I0�U�E�B@�H���M��]��E�M�@0�IP�U�E�BH�H8���M��]�E�M�@H�I �U�E�B�HP���M��]��E�M�@�I8�U�E�B0�H ���M��]��   �u��}�E_^[��]������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���   SVW�M��M��i���M����i���M���0�zi���M���H�oi�������$�����$�����$��\�����X���M����P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$��t����X���M������P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�M��EX���M���0���P�Q�P�Q�P�Q�P�Q�@�A�����$�����$�����$�M���W���M���H���P�Q�P�Q�P�Q�P�Q�@�A�E�_^[��]��������������������������������������������������������������������������������������������U���DSVW�M��EP�M��7U���EP�M����(U���EP�M���0�U���EP�M���H�
U���E�_^[��]� �������������������������������U���DSVW�M��E�_^[��]� ��������U���\SVW�M��EP�M�Q�U�R�TZ	�Hh�Q,�҃��M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[��]� �����������������������U���\SVW�M��EP�M�Q�U�R�TZ	�Hh�Q0�҃��M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[��]� �����������������������U���\SVW�M��EP�M�Q�U�R�TZ	�Hh�Q8�҃��M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[��]� �����������������������U���DSVW�M�_^[��]� �����������U����   SVW�M��}t
�   �B  �M���e���EP�M���M��Bx�ЉE؃}� u
�   �  �EP�M�=T���EԋM�9R���E�j/�E�P��Y����j�E�P��Y�����E�P�MQ�M�[[���E�    �	�E���E�}���   �}� uj �E�P�M��H���j �E�P�M��H���E�    �	�E����E��E�;E�}l�E�3�;E���;M�t�ݍ�H����EY����H���P�M�Q�UR�E���M��B|�Ѓ}��u��H����*V���j j��H���P�M�cg����H����
V����>����   _^[��]� ������������������������������������������������������������������������������������������������������U���   SVW�M��M�� d���M�����c���M���0��c�������$��t�����T���E���t������x����P��|����H�U��P�M��H�U��P�����$�M��T���E����M���U��P�M��H�U��P�M��H�U��P�����$�M��KT���E���0�M���U��P�M��H�U��P�M��H�U��P�E��H��XH�E��@P    �E�_^[��]��������������������������������������������������������������������������������U���DSVW�M�_^[��]��������������U���DSVW�M��EP�M�Q�TZ	�BH��   �у�_^[��]� ���������������U���DSVW�M��E�P�TZ	�Qd�B<�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�U�R�TZ	�Hd�Q�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�U�R�TZ	�Hd�Qp�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Qd���   �Ѓ�_^[��]� �����������������������U���DSVW�M��   _^[��]� ������U���DSVW�M�_^[��]� �����������U���DSVW�M�_^[��]�$ �����������U���DSVW�M�3�_^[��]� ���������U���  SVW�M�j�EP�@Q������t�����   �E�P�M�f���E������E�    �	�E����E��EP�M���M��Bx��9E���   ��<�����T����<���P�M�Q�UR�E���M��B|�Ѓ}��u��<����Q��룋EP�MQ�U�R��<���P������Q�F����P�M�W����t%�E��E�j�EP�xP������u��<����[Q�����<����NQ���?����E�_^[��]� ������������������������������������������������������������������������������U���@SVW�E#E_^[��]�����������U���   SVW�M���\���P�TZ	�QH�M��B,�й   ���}�E_^[��]� �����������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Qd�B�Ѓ�_^[��]� ��������������������������U���|  SVW�M��M�h��P������P�M�P��P�M�Q�G������D�����R��j �M��i����������D���P�MQ�UR��������������B|�Ѝ�D���P�MQ�U�R�EP������Q��D����;�����ԋ�
�H�J�H�J�H�J�H�J�@�B�MQ�UR�E���M����   ��ǅ ���   ��D����EO���� ���_^[��]� �����������������������������������������������������������������������U���   SVWj �M��9?���E�M�@�	�U��E�M�@0�I���U�E�BH�H���]��E�M�@ �	�U�B�E�M�@8�I���U�E�BP�H���]��E�M�@(�	�U�B�E�M�@@�I���U�E�BX�H���]��E�M�@�I�U�E�B0�H ���M�U�AH�J(���]��E�M�@ �I�U�E�B8�H ���M�U�AP�J(���]��E�M�@(�I�U�E�B@�H ���M�U�AX�J(���]ȋE�M�@�I0�U�E�B0�H8���M�U�AH�J@���]ЋE�M�@ �I0�U�E�B8�H8���M�U�AP�J@���]؋E�M�@(�I0�U�E�B@�H8���M�U�AX�J@���]��E�M�@�IH�U�E�B0�HP���M�U�AH�JX���]�E�M�@ �IH�U�E�B8�HP���M�U�AP�JX���]��E�M�@(�IH�U�E�B@�HP���M�U�AX�JX���]��   �u��}�E_^[��]��������������������������������������������������������������������������������������������������������������������������������������������������U���DSVW�M��EP�M�Q�TZ	�B@�H8�у�_^[��]� ������������������U���DSVW�M��TZ	�PH�M��B$��_^[��]��������������U���   SVW�M���\���P�TZ	�QH�M��B<�й   ���}�E_^[��]� �����������������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�3�_^[��]� ���������U���DSVW�M��   _^[��]�$ ������U���DSVW�M�_^[��]� �����������U���DSVW�M�_^[��]� �����������U���DSVW�M�_^[��]� �����������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�3�_^[��]� ���������U���`  SVW�M�S`����tj �EP�MQ�7������u3��   j h   ������P�Z����j �EP�M Q�UR�EP������Q�  ���E�H��E��t�E�^��E�� t�E�c��E%�   t�E�6��E��t�E�1�h   ������P�MQ�URj�>N����_^[��]�����������������������������������������������������������U���DSVW�M��M��c�������_^[��]����������������U���DSVW�M��TZ	�P�M��B<��_^[��]��������������U���@SVW�EP�MQ�UR�EP�MQ�UR�^�����E�M���   �Eǀ�   7��Eǀ�   ���Eǀ�   ���Eǀ�   F��Eǀ�   h��Eǀ�   ���Eǀ�   @��Eǀ�   ��_^[��]��������������������������������������������̋�`L����������̋�`\����������̋�`l����������̋�`P����������̋�``����������̋�`p����������̋�`D����������̋�`T����������̋�`d����������̋�`t����������̋�`H����������̋�`X����������̋�`h�����������U���@SVW�E�8 t�E�Q�TZ	�B��у��E�     _^[��]��������������������������U���@SVWhﾭޡTZ	�H��@  �҃�_^[��]�������������������������U���@SVW�} t�EP�TZ	�Q��@  �Ѓ�_^[��]�������������������U���@SVW�EP�MQ�TZ	�B���  �у�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B��  �у�_^[��]���������������������U���@SVW�TZ	�H��   ��_^[��]�����������������U���@SVW�} t�E�x��u�   �3�_^[��]�������������������������U���DSVW�=TZ	 t3�}s	�E�   ��E�E�j j �M�Q�TZ	�B���   �у��j�EP�    ��_^[��]�����������������������U���DSVW�}s�E   �E��P�,>�����E��}� u3��:�} t�E��Pj �M�Q��9�����E�� �����E����E��XZ	   �E�_^[��]������������������������������U���DSVW�=TZ	 t3�}s	�E�   ��E�E�j j �M�Q�TZ	�B���   �у��j�EP� �����_^[��]�����������������������U���DSVW�=TZ	 t3�}s	�E�   ��E�E�j j �M�Q�TZ	�B���   �у��j�EP������_^[��]�����������������������U���DSVW�=TZ	 t3�}s	�E�   ��E�E�j j �M�Q�TZ	�B���   �у��j�EP�@�����_^[��]�����������������������U���DSVW�} t=�E�E��=XZ	 t�E�x��u�E��P�hZ������E�P�TZ	�Q��Ѓ�_^[��]������������������������������U���DSVW�} t=�E�E��=XZ	 t�E�x��u�E��P��Y������E�P�TZ	�Q��Ѓ�_^[��]������������������������������U���@SVW�EP�TZ	�Q��Ѓ�_^[��]�������������U���@SVW�EP�TZ	�Q��Ѓ�_^[��]�������������U���DSVW�=TZ	 t7�}s	�E�   ��E�E��MQ�UR�E�P�TZ	�Q���   �Ѓ��j�EP������_^[��]�����������������������������������U���DSVW�=TZ	 tv�} t9�}s	�E�   ��E�E��MQ�UR�E�P�TZ	�Q���   �Ѓ��I�7�}s	�E�   ��E�E��MQ�UR�E�P�TZ	�Q���  �Ѓ���EP�MQ�������_^[��]��������������������������������������������������U���HSVW�} w�E   �=TZ	 t$�EP�MQ�UR�TZ	�H���   �҃��E��j�EP�B������E��M��M��E���thX���@	��
P�1�����E�_^[��]�����������������������������������������������U���@SVW�EP�MQ�TZ	�B��0  �у�_^[��]���������������������U���HSVW�} w�E   �=TZ	 tT�} t$�EP�MQ�UR�TZ	�H���   �҃��E��"�EP�MQ�UR�TZ	�H���  �҃��E��E��E��j�EP�"������E��E���thX���@	��P�0�����E�_^[��]�����������������������������������������������������U���@SVW�EP�TZ	�Q��Ѓ�_^[��]�������������U���@SVW�EP�TZ	�Q��Ѓ�_^[��]�������������U���@SVW�EP�TZ	�Q��Ѓ�_^[��]�������������U���@SVW�EP�TZ	�Q��Ѓ�_^[��]�������������U���@SVW�TZ	�H���   ��_^[��]�����������������U���@SVW�E�Q�TZ	�B���   �у��E�     _^[��]��������������U���DSVW�M��E�P�TZ	�Q���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�B���   �у�_^[��]� ���������������U���@SVW�TZ	�H���_^[��]���������������������U���@SVW�E�Q�TZ	�B�H�у��E�     _^[��]�����������������U���@SVW�E�Q�TZ	�B�H�у��E�     _^[��]�����������������U���XSVW�M�h�  �E�P�M�Q�TZ	�B���   �у�����V���E��M��9R���E�_^[��]������������������������U���DSVW�M��E�P�TZ	���   ��Ѓ�_^[��]�����������������������U���DSVW�M��E�P�TZ	���   �B8�Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�Q�B�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�B�H\�у�_^[��]� ������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�H���   �҃�_^[��]� ����������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�B�HX�у�_^[��]� ����������������������U���DSVW�M��E�P�TZ	�Q�B �Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�B���   �у�_^[��]� �������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q�B�Ѓ�_^[��]� ��������������������������U���@SVW�EP�MQ�UR�EP�MQ�TZ	�B��   �у�_^[��]�������������������������U���DSVW�M��EP�MQ�UR�EP�TZ	�Q�M��B$��_^[��]� ��������������������������U���DSVW�M��EP�MQ�TZ	�B�M���x  ��_^[��]� ���������������U���DSVW�M��TZ	�P�M���|  ��_^[��]�����������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�B�H(�у�_^[��]� ����������������������U���DSVW�M��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P�TZ	�Q�B`�Ѓ�(_^[��]�$ ����������������������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�B�H,�у�_^[��]� ����������������������U���DSVW�M��EP�MQ�UR�M��O����P�M���R����Pj j �E�P�TZ	�Q�B4�Ѓ� _^[��]� ������������������������������U���DSVW�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�TZ	�B�H4�у� _^[��]� ��������������������������U���DSVW�M��EP�MQ�U�R�TZ	�H�Q@�҃�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�B�HD�у�_^[��]� ������������������U���DSVW�M��E�P�TZ	�Q�BL�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�Q�BL�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�Q�BP�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�B�HT�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�B�HT�у�_^[��]� ������������������U���DSVW�M��EP�MQ�U�R�TZ	�H���   �҃�_^[��]� ����������������������������U���TSVW�M��EP�MQ�U�R�E�P�TZ	�Q���   �Ѓ�P�M�@���M��WJ���E_^[��]� �������������������U���DSVW�M��E��     �E��@    j �EP�M�Q�TZ	���   �H�у��E�_^[��]� �����������������������U���DSVW�M��E�P�TZ	�Q�Bh�Ѓ�_^[��]�������������������������U���HSVWh���@	��PhH_	h�   �[G�����E��}� t�M���L���E���E�    �E�_^[��]���������������������������������U���LSVW�E�8 t*�E��M��U��U��}� tj�M��J���E���E�    �E�     _^[��]����������������������U���DSVW�M��M��-���E��t�E�P�)�����E�_^[��]� ����������������������������U���DSVW�M��M�����6���M���B���E�_^[��]������������������������U���HSVW�M��M���E���E�    �	�E����E��}�}�E��M��D�    ��E�_^[��]���������������������������U���DSVW�M��M��5���M����1��_^[��]�����������U���DSVW�M��M���)��_^[��]����������������������U���DSVW�M��E��     �E��@`    �E��@d    �E��@h    �E����Xp�E��@x�����E��@|   _^[��]���������������������������U���DSVW�M��E��8 t j j j�E���P�M��	��C���E��     �E��x` t�E���`P�!����_^[��]������������������������������U���DSVW�M��E��8 th���@	��P�Z!�����E��x` th���@	��P�;!�����M��14���M���@���E�P�M���dQ�U��BxP�MQ�U���`R�dE�����M��A|�E��x|u�E��8 u>�E��8 u�E��x|u
�E��@|�����E��     �E���`P�� �����E��@|�   �E��xd ��   �E���pP�M���hQ�UR�9������u(�E��@h    �E����Xph���@	��P�^ �����EP�M����E��j j j�E���P�M��	�1B���U��B|�E��x|t�M��3���E��@|��E��@x�����E��@|_^[��]� ������������������������������������������������������������������������������������������������������������U���DSVW�M��M��~2���M��-?��_^[��]��������������U���DSVW�M��E��xd u�E��@`�}�E��M;Hxu�E��@`�j�EP�M��Q`Rj�E���P�M��	�A���U��B|�E��x|u �E��M�Hx�} t	�E�    �E��@`��E��@x�����} t�E�M��Q|�3�_^[��]� ���������������������������������������������U���DSVW�M��} t�E�M��Ap��E��xd t�E��@h��E��x|u�   �3�_^[��]� �����������������������U���@SVW�TZ	�H���_^[��]���������������������U���@SVW�E�Q�TZ	�B�H�у��E�     _^[��]�����������������U���DSVW�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�TZ	�B�H�у� _^[��]� ��������������������������U���DSVW�M��EP�M�Q�TZ	�B�H�у�_^[��]� ������������������U���DSVW�M��E�P�TZ	�Q�B�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�U�R�TZ	�H�Q�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�M��u�����M��k���H �F@��_^[��]� ���������������������U���DSVW�M��EP�MQ�UR�M��%�����M�����H �FD��_^[��]� ���������������������U���DSVW�M��M������xH u3���M��������M������H �FH��_^[��]������������������U���DSVW�M��M�����xL u3��&�EP�MQ�UR�M��s�����M��i���H �FL��_^[��]� �������������������U���DSVW�M��M��1���xP u����*�EP�MQ�UR�EP�M�������M�����H �VP��_^[��]� ������������������������������U���DSVW�M��M������xT u����"�EP�MQ�M�������M�����H �VT��_^[��]� ����������������������U���DSVW�M��M��a���xX u�����EP�M��J�����M��@���H �VX��_^[��]� ��������������������������U���lSVW�M��} t3�M������E�P�M��������M������H �VL�ҋM��M��h���} t9�M���:��P�M����M������M�����@@�E�}� t�E�P�M����_^[��]� �����������������������������������U���DSVW�M��E�P�MQ�TZ	�B�H�у��E�_^[��]� ���������������U���DSVW�M��M�����x` u� }  ��EP�M��������M������H �V`��_^[��]� ������������������������U���DSVW�M��EP�M�������M�����H �VH��_^[��]� �������������U���HSVW�M�j�EP�>���������P�M��u���E��M� C��;E��M�?��;E�~������*�EP�MQ�UR�EP�M�� �����M�����H �VD��_^[��]� ��������������������������������U���@SVW�E#E_^[��]�����������U���DSVW�M��M�����xP u������2�EP�MQ�UR�EP�MQ�UR�M�������M��z���H �FP��_^[��]� ������������������������������������U���DSVW�M��M��1���xT u������"�EP�MQ�M�������M��
���H �VT��_^[��]� ��������������������U���DSVW�M��M������xX u��EP�M�������M�����H �VX��_^[��]� �����������������������������U���XSVW�M��,���E�P�MQ�Y?������t�}� u3���E�P�M�Q�U�R�E�P�M���5��_^[��]�����������������������������������U���DSVW�M��E��     �E��@    �M��A    �U��B    �E��@    �E��@    �E�_^[��]��������������������������������U���PSVW�M��M�L9���M��-#����uh���@	��P�~����3��   �E�    �E�P�M�Q�UR�E�P�TZ	�Q���   �Ѓ���u3��M�E�    �	�E����E��E�;E�}"�E��M�<� u��E��M��R�M�;'���͍E�P�E&�����   _^[��]� ����������������������������������������������������������U���TSVW�M��M����M��-"����uh���@	��P�~����3��   �E�    �E�P�M�Q�UR�E�P�TZ	�Q���   �Ѓ���u3��o�}� u3��e�E�    �	�E����E��E�;E�}:�E��M�<� t�E��M���!����u�ϋE��M���U��E�P�M���뵍E�P�#%�����   _^[��]� ������������������������������������������������������������������������U���@SVW�TZ	�H��   ��_^[��]�����������������U���@SVW�E�Q�TZ	�B��$  �у��E�     _^[��]��������������U���DSVW�M��E�P�MQ�TZ	�B��(  �у��E�_^[��]� ����������������������������U���DSVW�M��E�P�MQ�TZ	�B��,  �у�_^[��]� ���������������U���DSVW�M��E�P�MQ�TZ	�B��,  �у������_^[��]� ������������������������U���@SVW�TZ	�H��0  ��_^[��]�����������������U���@SVW�TZ	�H��4  ��_^[��]�����������������U���@SVW�TZ	�H��p  ��_^[��]�����������������U���@SVW�TZ	�H��t  ��_^[��]�����������������U���HSVW�M��} t�M�('���E���E�    �E�P�M�Q�TZ	�B��8  �у�_^[��]� ���������������������U���DSVW�M��E��@_^[��]��������U���DSVW�M��EP�M�Q�TZ	�B��<  �у�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q��@  �Ѓ�_^[��]� �����������������������U���DSVW�M��EP�MQ�U�R�TZ	�H��D  �҃�_^[��]� ����������������������������U���DSVW�M��EP�M�Q�TZ	�B��H  �у�_^[��]� ���������������U���TSVW�M��EP�M�Q�U�R�TZ	�H��L  �҃�P�M�s4���M�����E_^[��]� ������������������������U���DSVW�M��E�P�TZ	�Q��T  �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�B��l  �у�_^[��]� ���������������U���DSVW�M��E�P�TZ	�Q��P  �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�B��X  �у�_^[��]� ���������������U���@SVW�TZ	�H��\  ��_^[��]�����������������U���@SVW�E�Q�TZ	�B��`  �у��E�     _^[��]��������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�H��d  �҃�_^[��]� ����������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�H��h  �҃�_^[��]� ����������������U���HSVW�M��E��8 t�E��H���M��	�E����E��}� |��E��@    _^[��]�����������������������������U���LSVW�M�j�M��q���E��EP�M�Q�m�����E�3�t�E��H���U��J�E�_^[��]� ���������������������U���HSVW�M��E��8 t�E��H���M��	�E����E��}� |��E��@    _^[��]�����������������������������U���LSVW�M�j�M��9+��Pj��7�����E��}� t�EP�m*�����M����E��E���E�    �E�_^[��]� ������������������������U���@SVW�E_^[��]��������������U���TSVW�M��E��HM�M��E��H�U�����M�E��M�;H��   j�EP�M��QR��6�����E�E�P�M���Q�U��P�M�����P�-�����E�}� tW�E��u-�E��8 t%�E��HQ�U�R�E��Q�u�����E�P������E��M��E��M�H�E��H�U���E��	�E��H�M��E��M��H�E�_^[��]� ����������������������������������������������������������������U���HSVW�EEk��+����E��E���}�U��}� u�}� u�E+E�E��E��E�_^[��]���������������������������U���TSVW�M��E��HM�M��E��H�U�����M�E��M�;H��   j�EP�M��QR�L5�����E�E�P�M���Q�U��P�M��~��P�?'�����E�}� tW�E��u-�E��8 t%�E��HQ�U�R�E��Q�u�����E�P�L�����E��M��E��M�H�E��H�U���E��	�E��H�M��E��M��H�E�_^[��]� ����������������������������������������������������������������U���HSVW�EPj�4�����E��}� t�M��U���M��M���E�    �E�_^[��]������������������������������U���DSVW�M��E�_^[��]�����������U���DSVW�M��E�_^[��]�����������U���@SVW�E��P�MQ�UR�E����_^[��]����������U���HSVW�E� h�   h@��M��T��P�EP�MQ������_^[��]������������������������U���DSVW�M��E��M��E��M�H�E�_^[��]� �����������������������U���@SVW�M���P�M�4��P�EP�MQ�TZ	�B��  �у�_^[��]�������������������U���DSVW�M��E�� _^[��]���������U���DSVW�M��E��@%��� _^[��]�������������������U���@SVW�E��P�MQ�UR������_^[��]����������U���HSVW�E� h�   h@��M�����P�EP�MQ�����_^[��]������������������������U���@SVW�E_^[��]��������������U���DSVW�E��M��E�P������E�     _^[��]��������������������U���DSVW�E��M��E�P�@�����E�     _^[��]��������������������U���DSVW�M��M��&���E�P�TZ	�Q$�BD�Ѓ��E�_^[��]��������������U���DSVW�M��M��u&���E�P�TZ	�Q$�BD�Ѓ��EP�M�Q�TZ	�B$�Hd�у��E�_^[��]� ����������������������������������U���DSVW�M��M��&���E�P�TZ	�Q$�BD�Ѓ��EP�M�Q�TZ	�B$�H�у��E�_^[��]� ����������������������������������U���DSVW�M��M��%���E�P�TZ	�Q$�BD�Ѓ��E�P�MQ�TZ	�B$�HL�у��E�_^[��]� ����������������������������������U���DSVW�M��E�P�TZ	�Q$�BH�Ѓ��M��<��_^[��]�����������������U���DSVW�M��EP�M�Q�TZ	�B$�HL�у�_^[��]� ������������������U���DSVW�M��EP�MQ�UR�EP�TZ	�Q$�M��B��_^[��]� ��������������������������U���DSVW�M��EP�TZ	�Q$�M��Bl��_^[��]� ����������������������U���DSVW�M��TZ	�P$�M��Bp��_^[��]��������������U���DSVW�M��E�P�TZ	�Q$�B�Ѓ�_^[��]�������������������������U���TSVW�M��E�P�M�Q�TZ	�B$�H�у�P�M�i'���M�����E_^[��]� ������������������������������U���DSVW�M��EP�M�Q�TZ	�B$�H�у�_^[��]� ������������������U���`SVW�M��E�P�M�Q�TZ	�B$�H �у�P�M�2'���M��\	���E_^[��]� ������������������������������U���`SVW�M��E�P�M�Q�TZ	�B$�H$�у�P�M��&���M������E_^[��]� ������������������������������U���`SVW�M��EP�M�Q�M��O����� ���M�����E_^[��]� �������������������������U���DSVW�M��E�P�TZ	�Q$�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�Q$�Bh�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�B$�H,�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�B$�H0�у�_^[��]� ������������������U���TSVW�M��E�P�M�Q�TZ	�B$�Ht�у�P�M�$���M�������E_^[��]� ������������������������������U���DSVW�M��EP�M�Q�TZ	�B$�H4�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�B$�H8�у�_^[��]� ������������������U���DSVW�M��E�P�MQ�TZ	�B$�HL�у��E�_^[��]� ���������������U���\SVW�EP�M��$���EP�M�Q�TZ	�B$�H@�у��E�P�M��#���M�� ���E_^[��]���������������������U���DSVW�M��EP�M�Q�TZ	�B$�H@�у��E�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�B$�H<�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�B$�H<�у������_^[��]� ���������������������������U���DSVW�M��EP�MQ�U�R�TZ	�H$�QP�҃�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�B$�HT�у�_^[��]� ������������������U���@SVW�TZ	�H$�QX��_^[��]��������������������U���@SVW�EP�TZ	�Q$�B\�Ѓ�_^[��]������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q$�B`�Ѓ�_^[��]� ��������������������������U���@SVW�TZ	�H(���_^[��]���������������������U���@SVW�E�Q�TZ	�B(�H�у��E�     _^[��]�����������������U���DSVW�M��EP�MQ�UR�EP�MQ�UR�TZ	�P(�M��B��_^[��]� �������������������U���DSVW�M��TZ	�P(�M��B��_^[��]��������������U���DSVW�M��EP�TZ	�Q(�M��B��_^[��]� ����������������������U���DSVW�M��EP�MQ�UR�TZ	�P(�M��B��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�B(�M��P ��_^[��]� ������������������U���DSVW�M�j�EP�MQ�TZ	�B(�M��P��_^[��]� ����������������U���DSVW�M��EP�MQ�UR�TZ	�P(�M��B$��_^[��]� ���������������U���DSVW�M��TZ	�P(�M��B(��_^[��]��������������U���DSVW�M��TZ	�P(�M��B,��_^[��]��������������U���DSVW�M��TZ	�P(�M��B0��_^[��]��������������U���DSVW�M��EP�TZ	�Q(�M��B4��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M��BX��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M��B\��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M��B`��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M��Bd��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M��Bh��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M��Bl��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M��Bx��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q(�M��Bt��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q(�M��Bp��_^[��]� ����������������������U���HSVW�M��EP�M�������t/�M��Q�M�������t�U��R�M������t	�E�   ��E�    �E�_^[��]� ����������������������������������U���HSVW�M��EQ� �$�M������t5�MQ�A�$�M�������t�UQ�B�$�M�������t	�E�   ��E�    �E�_^[��]� ���������������������������������������U���HSVW�M��EP�M������t/�M��Q�M������t�U��R�M������t	�E�   ��E�    �E�_^[��]� ����������������������������������U���HSVW�M��E��� �$�M��m�����t9�M���A�$�M��U�����t!�U���B�$�M��=�����t	�E�   ��E�    �E�_^[��]� ���������������������������������U���HSVW�M��EP�M��	����tB�M��Q�M��	����t/�U��R�M��v	����t�E��$P�M��c	����t	�E�   ��E�    �E�_^[��]� �������������������������������U���HSVW�M��EP�M�������tB�M��Q�M������t/�U��R�M������t�E��$P�M������t	�E�   ��E�    �E�_^[��]� �������������������������������U���HSVW�M��EP�M��c�����tB�M��Q�M��P�����t/�U��0R�M��=�����t�E��HP�M��*�����t	�E�   ��E�    �E�_^[��]� �������������������������������U���HSVW�M��EP�M������tB�M��Q�M��{����t/�U��0R�M��h����t�E��HP�M��U����t	�E�   ��E�    �E�_^[��]� �������������������������������U���\SVW�M��E�    �E�    �E�P�M��z�����u3��   �}� u#�M��j��P�M�����M������   �   h���@	��P�M�Q�TZ	�B���   �у��E�}� uj��M�����3��Lj �E�P�M�Q�M��	�����u�E�P�D����3��&j �E���P�M�Q�M�w���E�P������   _^[��]� ��������������������������������������������������������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q�B�Ѓ�_^[��]� ��������������������������U���\SVW�M��M�����E�P�M��;����u�E�    �M��"����E���E�P�M�]����E�   �M������E�_^[��]� ���������������������������������U���HSVW�M��E�P�M�������u3���E�����؋M��   _^[��]� �������������������U���DSVW�M��} ����Q�M�����_^[��]� ������������������������U���TSVW�M�j �M� �����E�h���@	��P�M�Q�TZ	�B���   �у��E��}� uj��M����3��[j �E�P�M�Q�M����E�P�M��b�����t�M�Q�U�R�M�������t	�E�   ��E�    �E��E��E�P� �����E�_^[��]� ���������������������������������������������������U���DSVW�M��EP�TZ	�Q�M��Bd��_^[��]� ����������������������U���DSVW�M��EP�MQ�UR�TZ	�P�M��Bh��_^[��]� ���������������U���XSVW�M��E�P�M�r���P�M�����E��M������E�_^[��]� ������������������������U���DSVW�M��EP�TZ	�Q(�M��B8��_^[��]� ���������������������U���DSVW�M��EP�TZ	�Q(�M��B<��_^[��]� ���������������������U���DSVW�M��EP�TZ	�Q(�M��B@��_^[��]� ���������������������U���DSVW�M��EP�TZ	�Q(�M��BD��_^[��]� ���������������������U���DSVW�M��EP�TZ	�Q(�M��BH��_^[��]� ����������������������U���DSVW�M��EP�MQ�TZ	�B(�M��P|��_^[��]� ������������������U���DSVW�M��EP�TZ	�Q(�M��BL��_^[��]� ����������������������U���DSVW�M��EP�MQ�TZ	�B(�M����   ��_^[��]� ���������������U���DSVW�M����E�$�TZ	�P(�M��BT��_^[��]� ������������������U���DSVW�M�Q�E�$�TZ	�P(�M��BP��_^[��]� ��������������������U���@SVW�TZ	�H(�Q��_^[��]��������������������U���@SVW�E�Q�TZ	�B(�H�у��E�     _^[��]�����������������U���DSVW�M��E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP�TZ	�Q(�M����   ��_^[��]�( �������������������������������U���@SVW�EP�MQ�UR�EP�MQ�TZ	�B(�H�у�_^[��]����������������������������U���@SVW�TZ	�H,�Q,��_^[��]��������������������U���DSVW�M��TZ	�P,�M��B4��_^[��]��������������U���@SVW�E�Q�TZ	�B,�H0�у��E�     _^[��]�����������������U���DSVW�M��TZ	�P,�M��B8��_^[��]��������������U���`SVW�M��E�P�TZ	�Q,�M��B<��P�M�����M�� ����E_^[��]� ������������������U���TSVW�M��EP�M�Q�TZ	�B,�M��P@��P�M�9���M������E_^[��]� ������������������������������U���@SVWj j �TZ	�H,��҃�_^[��]��������������U���DSVW�M��EP�MQ�U�R�TZ	�H,�Q�҃�_^[��]� ���������������U���@SVW�E�Q�TZ	�B,�H�у��E�     _^[��]�����������������U���DSVW�M��TZ	�P,�M��B��_^[��]��������������U���DSVW�M��TZ	�P,�M��B��_^[��]��������������U���DSVW�M��TZ	�P,�M��B��_^[��]��������������U���DSVW�M��TZ	�P,�M��B ��_^[��]��������������U���DSVW�M��TZ	�P,�M��B$��_^[��]��������������U���DSVW�M��TZ	�P,�M��B(��_^[��]��������������U���DSVW�M��EP�MQ�TZ	�B,�M��P��_^[��]� ������������������U���`SVW�M��E�P�TZ	�Q,�M��B��P�M�6���M��`����E_^[��]� ������������������U���@SVW�EP�MQ�UR�TZ	�H��D  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H��H  �҃�_^[��]������������������U���@SVW�EP�TZ	�Q��L  �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�TZ	�B�H�у�_^[��]������������������������U���@SVW�EP�MQ�UR�TZ	�H�Q�҃�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B�H�у�_^[��]������������������������U���@SVW�EP�MQ�UR�TZ	�H�Q�҃�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B�H�у�_^[��]������������������������U���@SVW�EP�MQ�TZ	�B���  �у�_^[��]���������������������U���@SVW�EP�TZ	�Q�B�Ѓ�_^[��]������������U���lSVW�E�P�M�i����M��4�����u�E�    �M������E��~j�E�P�F�������u$�E�P�������u�E�    �M��l����E��Hj�EP��������u$�EP�>������u�E�    �M��6����E���E�   �M��"����E�_^[��]�������������������������������������������������������U���@SVW�EP�TZ	�Q�B �Ѓ�_^[��]������������U���@SVW�EP�MQ�TZ	�B�H(�у�_^[��]������������������������U���@SVW�EP�MQ�UR�EP�MQ�TZ	�B��  �у�_^[��]�������������������������U���@SVW�EP�MQ�UR�EP�TZ	�Q��   �Ѓ�_^[��]�����������������������������U���@SVW�EP�TZ	�Q��  �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�UR�TZ	�H��  �҃�_^[��]������������������U���\SVW�E�P�TZ	�Q�B$�Ѓ�P�M�����M��#����E_^[��]������������������������U���\SVW�E�P�TZ	�Q���  �Ѓ�P�M����M�������E_^[��]���������������������U���@SVW�EP�MQ�TZ	�B���  �у�_^[��]���������������������U���   SVW�E�    �=tZ	 t�E�P�tZ	������M���|�����M�����M���|�����|����M��U�R�M�����E���t�e���M�� ����M���t�e���M�������E_^[��]�������������������������������������������������U���\SVW�EP�M�Q�TZ	�B���  �у�P�M�R���M��|����E_^[��]�����������������U���@SVWj�EP��������E_^[��]����������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�TZ	�H���   ��_^[��]�����������������U���@SVW�EP�TZ	�Q���   �Ѓ��E�     _^[��]����������������U���DSVW�M��EP�MQ�UR�EP�TZ	�Q�M����_^[��]� ���������������������������U���DSVW�M��TZ	�P�M��B��_^[��]��������������U���DSVW�M��TZ	�P�M����   ��_^[��]�����������U���DSVW�M��EP�TZ	�Q�M��B`��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��Bd��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��Bh��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��Bl��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��Bp��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��Bt��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M���  ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M��Bx��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M��B|��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�M�Q�TZ	�B��  �у�_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�B�M����   ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�B�M����   ��_^[��]� ���������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���HSVW�M��} t&�EP�M�Q�TZ	�B �H$�у���t	�E�   ��E�    �E�_^[��]� ���������������������U���DSVW�M��E�P�MQ�UR�TZ	�H �QL�҃�_^[��]� ���������������U���DSVW�M��} u3���EP�M�Q�TZ	�B �H(�у��   _^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M��B��_^[��]� ���������������������U���DSVW�M��EP�TZ	�Q�M��B��_^[��]� ���������������������U���DSVW�M��EP�TZ	�Q�M��B��_^[��]� ���������������������U���DSVW�M��EP�TZ	�Q�M��B��_^[��]� ���������������������U���DSVW�M��EP�TZ	�Q�M��B��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��B��_^[��]� ����������������������U���DSVW�M��EP�MQ�TZ	�B�M��P\��_^[��]� ������������������U���DSVW�M��EP�MQ�TZ	�B�M���  ��_^[��]� ���������������U���DSVW�M����E�$�TZ	�P�M��B ��_^[��]� ������������������U���DSVW�M�Q�E�$�TZ	�P�M��B$��_^[��]� ��������������������U���DSVW�M����E�$�TZ	�P�M��B(��_^[��]� ������������������U���DSVW�M��EP�TZ	�Q�M��B,��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��B0��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��B4��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��B8��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��B<��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��B@��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��BD��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��BH��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��BL��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M��BP��_^[��]� ����������������������U���DSVW�M��EP�MQ�UR�EP�TZ	�Q�M����   ��_^[��]� �����������������������U���DSVW�M��EP�TZ	�Q�M��BT��_^[��]� ����������������������U���DSVW�M��EP�M�Q�TZ	�B��  �у�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�EP�TZ	�Q�M����   ��_^[��]� �����������������������U���DSVW�M��EP�MQ�UR�EP�TZ	�Q�M����   ��_^[��]� �����������������������U���DSVW�M��EP�MQ�TZ	�B�M��PX��_^[��]� ������������������U���DSVW�M��TZ	�P�M����   ��_^[��]�����������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���DSVW�M��EP�MQ�TZ	�B�M����   ��_^[��]� ���������������U���DSVW�M��TZ	�P�M����   ��_^[��]�����������U���DSVW�M��EP�MQ�TZ	�B�M����   ��_^[��]� ���������������U���DSVW�M��TZ	�P�M����   ��_^[��]�����������U���DSVW�M��TZ	�P�M����   ��_^[��]�����������U���DSVW�M��TZ	�P�M����   ��_^[��]�����������U���@SVW�EP�MQ�UR�EP�MQ�TZ	�B���   �у�_^[��]�������������������������U���@SVW�EP�MQ�UR�EP�TZ	�Q��   �Ѓ�_^[��]�����������������������������U���PSVW�EP�MQ�U�R�TZ	�H���  �҃�P�M�V����M������E_^[��]������������������������������U���@SVW�EP�MQ�TZ	�B���  �у�_^[��]���������������������U���PSVW�M��M�;����E��}�NIVbP�}�NIVb��   �}�TCAb,�}�TCAb�7  �}�$'  �j  �}�MicM��   �p  �}�INIbtJ�b  �}�atni$�}�atnit)�}�ckhc�  �}�ytsdtL�5  �}�cnyst�'  ������  �E��x t
�   �  �E��@   �E���M��B����   �E���M��B�ЋE��@    ��   �E��x u
�   ��   �E���M��B���   j hIicM�M�>����E��EP�M�Q�U���M��P���   j hIicM�M�����E��EP�M�Q�U���M��P���Zj hdiem�M������E��EP�M�Q�U���M��P�҉E�E��+�E���M��B�����EP�M���M��B�и   �3�_^[��]� �����������������������������������������������������������������������������������������������������������������������������������U���DSVW�M��TZ	�P�M��B ��_^[��]��������������U���DSVW�M��E�� l��E�Ph��TZ	�Q0��Ѓ��M��A�E��@    �E�_^[��]�������������������������U���lSVW�E�    �M�������} tO�EP�TZ	�Q4�B�Ѓ��E�}� u�E�    �M��b����E��   �E�P�MQ�U��M�P(�҉E��J�EP�TZ	�Q0�B�Ѓ��E��}� u�E�    �M������E��O�E�P�MQ�U���M��P �҉E��M��������t�E�P�MQ�TZ	�B0�Hx�у��E��E��M�������E�_^[��]����������������������������������������������������������������������������U���DSVW�M��M�������E��t�E�P��������E�_^[��]� ����������������������������U���DSVW�M��E�� l��E��x t�E��HQ�TZ	�B0�H�у��E��@    _^[��]��������������������������U���DSVW�M��E��HQ�TZ	�B0���   �у�_^[��]�������������������U���DSVW�M��EP�M��QR�TZ	�H0���   �҃�_^[��]� �������������U���DSVW�M��M��n���P�TZ	�H0���   �҃�_^[��]������������������U���DSVW�M�j j j j j j j j j4�E��HQ�TZ	�B0���   �у�(_^[��]�����������������U���DSVW�M�j j j j j j j j j;�E��HQ�TZ	�B0���   �у�(_^[��]�����������������U���DSVW�M��EP�M�����P�TZ	�Q0���   �Ѓ�_^[��]� ��������������������������U���`SVW�M��E P�M������EPh8kds�M������E�    �E�P�M�Qj �UR�EP�MQ�UR�EPj2�M������P�TZ	�Q0���   �Ѓ�(�E�E��M������E�_^[��]� �����������������������������������������U���DSVW�M��M�����P�TZ	�H0���   �҃�_^[��]������������������U���DSVW�M��E��x u3��bj j j j j �E Pj �MQj�U��BP�TZ	�Q0���   �Ѓ�(�EP�MQ�UR�EPj �MQ�U��BP�TZ	�Q0���   �Ѓ�_^[��]� ��������������������������������������������U���DSVW�M��E��x u3���E��HQ�TZ	�B0�H�у�_^[��]�������������������������U���DSVW�M��M������_^[��]� �������������������U���TSVW�M��E��x uj �M�o����E�I�M�!���P�EP�M�{���P�M��QR�E�P�TZ	�Q0���   �Ѓ�P�M������M������E_^[��]� ������������������������������������������U���DSVW�M��E��    �E��M�H�E�_^[��]� ����������������������U���DSVW�M��E�� _^[��]���������U���DSVW�M��E��@_^[��]��������U���DSVW�M��EP�M��QR�TZ	�H0�Q�҃�_^[��]� ����������������U���DSVW�M��E��x u�.j j j j j j �EPj j�M��QR�TZ	�H0���   �҃�(_^[��]� ����������������������������������U���DSVW�M��E��x u3��-�M�\���P�EP�M����P�M��QR�TZ	�H0�Q�҃�_^[��]� ���������������������������������U���DSVW�M��E��x u3��-�M�����P�M�J���P�E��HQ�TZ	�B0���   �у�_^[��]� ���������������������������������U���DSVW�M��E��x u3��-�M�|���P�EP�M�����P�M��QR�TZ	�H0�Q\�҃�_^[��]� ���������������������������������U���DSVW�M��E��x u3��#�EP�MQ�U��BP�TZ	�Q4��  �Ѓ�_^[��]� ���������������������������U���DSVW�M��E��x u3�� �EP�MQ�U��BP�TZ	�Q4�Bh�Ѓ�_^[��]� ������������������������������U���DSVW�M��E��x u3�� �EP�MQ�U��BP�TZ	�Q4�Bp�Ѓ�_^[��]� ������������������������������U���DSVW�M��E��x u3��#�EP�MQ�U��BP�TZ	�Q4��  �Ѓ�_^[��]� ���������������������������U���DSVW�M�h���h  ��EPj 3Ƀ} ����Qj �UR�EP�M��i���_^[��]� ����������������������������U���lSVW�M�htniv�M��?����EPhulav�M������hgnlfhtmrf�M�������EPhinim�M�������EPhixam�M�������EPhpets�M������EPhsirt�M������}   �u	�}$���t"�E Ph2nim�M��{����E$Ph2xam�M��j����E�P�MQ�U�R�M��������J����E��M������M������E�_^[��]�  ������������������������������������������������������������������U���lSVW�M�htlfv�M��������E�$hulav�M�蹺���E,Phtmrf�M��������E�$hinim�M�蒺�����E�$hixam�M��|������E$�$hpets�M��f����EDPhsirt�M��[����E0��������Dz�E8��������D{,���E0�$h2nim�M��#������E8�$h2xam�M������E@Phdauq�M������E�P�MQ�U�R�M�������������E��M��6����M�裼���E�_^[��]�@ ��������������������������������������������������������������������������U���DSVW�M����E�$�EP�TZ	�Q�M��B,��_^[��]� �������������U���   SVW�M�hgnrs�M��\����EP��t���������t���Qj�M�褻����t����Q����EP�M������M�Qj�M������M��/����E�P�MQ�U�R�M��w����������E��M��	����M��v����E�_^[��]� ���������������������������������������������U���DSVW�M��E��    �E��M�H�E�_^[��]� ����������������������U���DSVW�M��EP�MQ�TZ	�B�M����   ��_^[��]� ���������������U���lSVW�M�hmnrs�M������EPj�M�������E�P�MQ�U�R�M��i����������E��M�������M��h����E�_^[��]� �������������������������������U���lSVW�M��E�����DSSSP�M�����j�M������P�M��7����E�P�MQ�U�R�M��پ���������E��M��k����M��ع���E�_^[��]� �������������������������������U���lSVW�M�hCITb�M�������EPhCITb�M��G����EPhsirt�M������EPhulav�M������E�P�MQ�U�R�M��4������r����E��M�������M��3����E�_^[��]� ������������������������������������������U���XSVW�M�j �EP�M�Q�M�,���P�UR�M��0����E��M��_����E�_^[��]� ������������������������������U���DSVW�M��E,Pj �����$�����$htemf���E$�$���E�$���E�$���E�$�MQ�M��m���_^[��]�( ��������������������������������U���TSVW�M��E���������Dz�E�]�����E�$�G������]��E���������Dz�E�]�����E�$�������]��E,Pj �����$�����$hrgdf���E$�$������$���E��$���E��$���E�$�MQ�M�����_^[��]�( ������������������������������������������������������������U���@SVW�E�ȴ�5��_^[��]������������������U���DSVW�M��E,Pj �����$�����$htcpf�E$�5H����$�E�5H����$�E�5H����$���E�$�MQ�M�����_^[��]�( ������������������������������U���DSVW�M��E��x u3��D�M����P�E P���E�$���E�$�MQ�M�����P�U��BP�TZ	�Q0�B(�Ѓ�$_^[��]� ��������������������������U���LSVW�M��E��x u3��A�M����P�E�P�M�v���P�M��QR�TZ	�H0�Q,�҃��E�3��}� ���M��E�_^[��]� �����������������������������U���DSVW�M��E��x u3��-�M����P�EP�M�����P�M��QR�TZ	�H0�Q,�҃�_^[��]� ���������������������������������U���DSVW�M��E��x u3��-�M�,���P�EP�M����P�M��QR�TZ	�H0�Q0�҃�_^[��]� ���������������������������������U���DSVW�M��EP�MQ�M�������u3��;�E��P�MQ�M��z�����u3�� �E��P�MQ�M��_�����u3���   _^[��]� ����������������������������������������U���XSVW�M��E��x u3��   �E�    �M�"���P�E�P�M�|���P�M��QR�TZ	�H0�Q8�҃��E�}� tG�}� tA�E�P�M�4����}� t(�E��E��M��M��}� tj�M��˱���E���E�    �E�    �E�_^[��]� ����������������������������������������������������U���DSVW�M��M�葱���E��t�E�P�j������E�_^[��]� ����������������������������U���`SVW�M��M������E�P�MQ�M�舴���E�}� u�E�    �M������E���E�P�M�T����E�E��M�������E�_^[��]� �������������������������U���DSVW�M��E��x u3��2�M�|���P�EP�MQ�M�����P�U��BP�TZ	�Q0�B<�Ѓ�_^[��]� ����������������������������U���LSVW�M��E�    �E�P�MQ�M��ݵ���E�E�P�MQ�M�����E�_^[��]� ������������������������������U���DSVW�M��EP�MQ�TZ	�B�M��P0��_^[��]� ������������������U���LSVW�M��E�P�MQ�M��{����E�E�P�MQ�M�/����E�_^[��]� ���������������������U���PSVW�M��E�P�MQ�M�������E����E��$�EP�M�ԭ���E�_^[��]� ����������������U���\SVW�M��M������E�P�MQ�M�������u3��E�E�P�MQ�M�������u3��-�E�P�MQ�M��m�����u3���E�P�MQ�M� ����   _^[��]� ��������������������������������������U���\SVW�M��M��E����E�P�MQ�M�踱���E�E�P�MQ�M�z����E�E��M��@����E�_^[��]� �������������������������������U���hSVW�M��M������E�P�MQ�M��a����E܍E�P�MQ�M�t����E܉E��M������E�_^[��]� �������������������������������U���DSVW�M��EP�MQ�TZ	�B�M��P<��_^[��]� ������������������U���hSVW�M��M�������E�P�M�Q�UR�M�萾���E؃}�t�E�P�MQ�M苹���}�t���E��$�EP�M蜫���E�_^[��]� ����������������������������������������U���DSVW�M�j j �EP�M�g���P�MQ�M�蚹��_^[��]� ��������������U���DSVW�M��EP�MQ�TZ	�B�M����   ��_^[��]� ���������������U���DSVW�M��E$P�M Qj �UR�EP�MQj �UR�M�b���P�EP�M������_^[��]�  ��������������������������U���DSVW�M�j �E@P���E8�$���E0�$�M,Q���E$�$���E�$���E�$�����$�UR�M�z������$�EP�M�����_^[��]�< ������������������������������U���DSVW�M����E�$�EP�TZ	�Q�M����   ��_^[��]� ��������������������������U���DSVW�M�j ���E$�$���E�$���E�$�����$�EP�M贿�����$�MQ�M�跹��_^[��]�$ ������������������������U���DSVW�M�j ���E$�$���E�$���E�$�����$�EP�M�D������$�MQ�M��~���_^[��]�$ ������������������������U���DSVW�M�j ���E$�$���E�$���E�$�����$�EP�M�Ծ�����$�MQ�M��g���_^[��]�$ ������������������������U���hSVW�M��EPj �M�����P�MQ�U�R�M�����P�EP�M��S����E��M�肩���M��z����E�_^[��]� �������������������������U���   SVW�M�j �M������P�EP�M�Q�M�*���P�UR�M�������E��M��`����M��X����E�_^[��]� ��������������������������U���`SVW�M��EP�MQ�U�R�TZ	�P�M����   ��P�M������M�������E_^[��]� ������������������������U���|SVW�M����]�}�t�����$�EP�M�6����]�E P���E�$���E��$�M�����P�MQ�U�R�M�����P�EP�M��f���_^[��]� �����������������������������U���xSVW�M��} u�TZ	�H���   �҉E�} u3��y  �M�����E�htlfv�M��~����M�����M����$�^������M�]��Q������$�E������}����$hulav�M������hmrffhtmrf�M������M謷���M����$�������M�]���������$��������}����$hinim�M�蜥���M�d����M����$�������M�]�诹�����$�������}����$hixam�M��T��������$hpets�M��?���j hdauq�M��6����E�Phspff�M��%����E Phsirt�M������E�P�MQ�U�R�M�趬����������E��M��H����M�赧���E�_^[��]� ����������������������������������������������������������������������������������������������������������������������������U���@SVW���E�$�7�����_^[��]����������������U���DSVW�M��E�� _^[��]���������U���DSVW�M��E��@_^[��]��������U���dSVW�M��} u�TZ	�H���   �҉E�} u3��`�M�p����E��E�P�MQ�M������E��E��ش���$�E��ش���$�M��`����M���P�Q�P�Q�@�A�E�_^[��]� ����������������������������������������U���dSVW�M�j �E P�MQ�UR�M��M���P�EP�M�Q�M�����P�UR�EP�M�����_^[��]� �������������������U���DSVW�M��E�����E����X�E�_^[��]������������U���TSVW�M��EP�MQ�U�R�TZ	�P�M����   �ЋM���P�Q�P�Q�@�A�E_^[��]� ��������������������������������U���XSVW�M��M��[����E�P�MQ�UR�M��u����E�E�P�MQ�M�
����E�_^[��]� �������������������������U���DSVW�M��EP�MQ�TZ	�B�M��P@��_^[��]� ������������������U���DSVW�M��E��x u3��;�M蜼��Pj j j j j j �M����Pj1�E��HQ�TZ	�B0���   �у�(_^[��]� �����������������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj j �MQ�UR�EP�MQ�URj�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���DSVW�M��E��x u3��.j j j j j j j �EPj-�M��QR�TZ	�H0���   �҃�(_^[��]� ��������������������������������U���HSVW�M��E��x u3��=�E�    �E�Pj j j �MQ�URj j j)�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������������U���HSVW�M��E��x u3��=�E�    �E�Pj j �MQj �URj j j)�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������������U���DSVW�M��E��x u3��4j j j �EP�MQ�URj �EPj/�M��QR�TZ	�H0���   �҃�(_^[��]� ��������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj j �MQ�UR�EP�MQ�URj'�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj j �MQ�UR�EP�MQ�URj,�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj j �MQ�UR�EP�MQ�URj�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��D�E�    �E�Pj �MQ�UR�EP�MQ�UR�EPj�M��QR�TZ	�H0���   �҃�(�E�_^[��]� ��������������������������U���DSVW�M�j j j �EP�MQ�URj �EPj.�M��QR�TZ	�H0���   �҃�(_^[��]� �����������������������U���HSVW�M��E��x u3��C�E�    �E�Pj �MQ�UR�EP�MQj �URj�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj �MQ�UR�EP�MQj �URj:�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj �MQ�UR�EP�MQj �URj�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj �MQ�UR�EP�MQj �URj*�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��A�E�    �E�Pj j �MQ�UR�EPj �MQj�U��BP�TZ	�Q0���   �Ѓ�(�E�_^[��]� �����������������������������U���HSVW�M��E��x u3��A�E�    �E�Pj j �MQ�UR�EPj �MQj�U��BP�TZ	�Q0���   �Ѓ�(�E�_^[��]� �����������������������������U���HSVW�M��E��x u3��A�E�    �E�Pj j �MQ�UR�EPj �MQj	�U��BP�TZ	�Q0���   �Ѓ�(�E�_^[��]� �����������������������������U���HSVW�M��E��x u3��A�E�    �E�Pj j �MQ�UR�EPj �MQj
�U��BP�TZ	�Q0���   �Ѓ�(�E�_^[��]� �����������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj �MQ�UR�EP�MQj �URj�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj �MQ�UR�EP�MQj �URj�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���DSVW�M��E��x u3��4j j j �EP�MQ�URj �EPj�M��QR�TZ	�H0���   �҃�(_^[��]� ��������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj �MQ�UR�EP�MQj �URj�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��C�E�    �E�Pj �MQ�UR�EP�MQj �URj>�E��HQ�TZ	�B0���   �у�(�E�_^[��]� ���������������������������U���HSVW�M��E��x u3��A�E�    �E�Pj j �MQ�UR�EPj �MQj�U��BP�TZ	�Q0���   �Ѓ�(�E�_^[��]� �����������������������������U���DSVW�M��E��x u3��?�M�l���Pj j j j �EP�MQ�M躨��Pj�U��BP�TZ	�Q0���   �Ѓ�(_^[��]� �������������������������������U���TSVW�M��EP�M��i����E�P�M�Q�M��ϱ����t+�}� u��M������P�E�P�MQ�M�蓹����u3�����   _^[��]� ���������������������������U���DSVW�M��E��x u3��;�M�l���Pj j j j j j �M辧��Pj�E��HQ�TZ	�B0���   �у�(_^[��]� �����������������������������������U���HSVW�M��E��x u3��A�E�    �E�Pj j �MQ�UR�EPj �MQj�U��BP�TZ	�Q0���   �Ѓ�(�E�_^[��]� �����������������������������U���DSVW�M��E��x u3��$�EP�MQ�UR�E��HQ�TZ	�B0�HD�у�_^[��]� ��������������������������U���DSVW�M��E��x u3��;�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U��BP�TZ	�Q0���   �Ѓ�$_^[��]�  �����������������������������������U���DSVW�M��E��x u3���E��HQ�TZ	�B0�HX�у�_^[��]�������������������������U���DSVW�M��E��x u3�� �EP�MQ�U��BP�TZ	�Q0�BL�Ѓ�_^[��]� ������������������������������U���DSVW�M��E��x u3�� �E   �P�M��QR�TZ	�H0�QP�҃�_^[��]� ������������������������������U���DSVW�M��E��x u3���EP�M��QR�TZ	�H0�QP�҃�_^[��]� �������������������U���DSVW�M��E��x u3��'�EP�MQ�UR�EP�M��QR�TZ	�H0�QT�҃�_^[��]� �����������������������U���DSVW�M��E�HQ�TZ	�B4��у��E�@    �E�M��H�M诫��P�EP�MQ�M����P�U��BP�TZ	�Q0���   �Ѓ��M�A�E3Ƀx ����_^[��]� ����������������������������������������U���DSVW�M��E��x u3��.j j j j j �EPj j j�M��QR�TZ	�H0���   �҃�(_^[��]� ��������������������������������U���DSVW�M��} u3��4�E�@    �M芧��P�EP�M��}���P�TZ	�Q0���   �Ѓ�_^[��]� �����������������������������U���DSVW�M�j j j j j j j j j0�M�����P�TZ	�H0���   �҃�(_^[��]��������������������������������U���DSVW�M��} u�E@Z	�EP�M�O���P�MQ�U��BP�TZ	�Q0�B@�Ѓ�_^[��]� ���������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U��BP�TZ	�Q0�Bd�Ѓ�_^[��]� �������������������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U��BP�TZ	�Q0�Bp�Ѓ�_^[��]� �������������������������������U���DSVW�M��M�ɨ��P�EP�MQ�UR�EP�M����P�M��QR�TZ	�H0�Qh�҃�_^[��]� ����������������������������������U���DSVW�M�j j j j j j j �M負��Pj�E��HQ�TZ	�B0���   �у�(_^[��]� �����������������������U���DSVW�M�j j j j j jj �M�R���Pj�E��HQ�TZ	�B0���   �у�(_^[��]� �����������������������U���DSVW�M�j j j j j j j �M����Pj�E��HQ�TZ	�B0���   �у�(_^[��]� �����������������������U���`SVW�M��M��(����M�1���P�E�Pj j j j j �M聟��Pj8�M��QR�TZ	�H0���   �҃�(�E�}� t�E�P�M�o����E�E��M��z����E�_^[��]� ���������������������������������U���DSVW�M��M虦��P�EPj j j j j �M����Pj9�M��QR�TZ	�H0���   �҃�(_^[��]� �������������������������������U���DSVW�M��M�)���Pj j j j j j �M�{���Pj"�E��HQ�TZ	�B0���   �у�(_^[��]� ��������������������������������U���DSVW�M��M蹥��Pj j j j j j �M����Pj5�E��HQ�TZ	�B0���   �у�(_^[��]� ��������������������������������U���DSVW�M��M�I���Pj j j j �EPj �M虝��Pj<�M��QR�TZ	�H0���   �҃�(_^[��]� �������������������������������U���DSVW�M�j j �EP�MQ�UR�EPj �MQj3�U��BP�TZ	�Q0���   �Ѓ�(_^[��]� ��������������������U���DSVW�M�j j j j j �EPj �MQj�U��BP�TZ	�Q0���   �Ѓ�(�EP�M��QR�TZ	�H0�Qt�҃�_^[��]� �������������������������������U���DSVW�M�j j j j j j �EPj j�M��QR�TZ	�H0���   �҃�(_^[��]� �����������������������������U���DSVW�M�j j j j j j j j j�E��HQ�TZ	�B0���   �у�(_^[��]�����������������U���DSVW�M�j j j j j j j �EPj�M��QR�TZ	�H0���   �҃�(_^[��]� �����������������������������U���DSVW�M�j j j j j j j j j(�E��HQ�TZ	�B0���   �у�(_^[��]�����������������U���DSVW�M�j j j j j j �EP�MQj&�U��BP�TZ	�Q0���   �Ѓ�(_^[��]� ��������������������������U���DSVW�M�j j j j �EP�MQj �URj+�E��HQ�TZ	�B0���   �у�(_^[��]� ������������������������U���DSVW�M�j j j j j j j j j�E��HQ�TZ	�B0���   �у�(_^[��]�����������������U���DSVW�M�j j j j j j j j j#�E��HQ�TZ	�B0���   �у�(_^[��]�����������������U���DSVW�M��} tj j�M褟���M��} tj j�M荟���M��EP�MQ�U��BP�TZ	�Q0�B`�Ѓ�_^[��]� �����������������������������U���DSVW�M��EP�MQ�UR�E��HQ�TZ	�B0���   �у�_^[��]� ��������������������U���DSVW�M�j j j j j j j j j �E��HQ�TZ	�B0���   �у�(_^[��]�����������������U���DSVW�M��   _^[��]���������U���DSVW�M��   _^[��]���������U���DSVW�M�_^[��]��������������U���DSVW�M��   _^[��]� ������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�3�_^[��]������������U���DSVW�M�_^[��]� �����������U���DSVW�M��M�辡���E�� ��E��@   �E��@    �E�_^[��]����������������������U���DSVW�M��M��W����E��t�E�P��������E�_^[��]� ����������������������������U���DSVW�M��E�� ��M�踞��_^[��]�������������U���HSVW�M��E��@    j �EP�MQ�UR�EPj 3Ƀ} ����
Q�M�������t�U��z t	�E�   ��E�    �E�_^[��]� ����������������������������������������U���DSVW�M��E��M�H�M��5���_^[��]� ����������U���PSVW�M��M������E��}�ckhc �}�ckhct,�}�cksatS�}�TCAbtf��   �}�atnit�   3��   �E��x t �M�������t�E��@    �   �   3��   �E��x t�E���M��B���t3��pj hdiem�M肛���E��E��@   �EP�M�Q�U���M��P�҉E�E��x t�}�t�}�u3��}���P�M�脬���E���EP�MQ�M�跑��_^[��]� ����������������������������������������������������������������������U���PSVW�M��E��x u��   �E�E��}���   �M��$��C�E;E~��   �   �E;E|�   �{�E;E}�   �l�E;E�   �]�E;E~�E;E}�   �F�E;E|
�E;E�v�2�E;E|
�E;E}�b��E;E~
�E;E�N�
�E;Et�B�EP�M������M�Q�M�耟��j�E���$�E���$�EP��������E��@    _^[��]� ��BCC$C3CJC^CrC�C��������������������������������������������������������������������������������U���DSVW�M��E��M��E��@    �E�_^[��]� ����������������������U���PSVW�M��E��x u�I  �E�E��}���   �M��$��E�E�]����z�  ��   �E�]����Az�  �   �E�]����Au��   �   �E�]����u��   �   �E�]����z�E �]����Au�   �n�E�]����Az�E �]����u�   �M�E�]����Az�E �]����Au�u�/�E�]����z�E �]����u�W��E�E������D{�D�EP�M������M�Q�M��a����E(P���E �$���E�$�MQ�ڂ�����E��@    _^[��]�$ �D�D�D	E EAEbE�E�E����������������������������������������������������������������������������������������������������������������U���DSVW�M�j���E �$���E�$���E�$�EP�MQ�M�蛃��_^[��]�  ������������������������������U���DSVW�M�j���E �$���E�$���E�$�EP�MQ�M��;���_^[��]�  ������������������������������U���DSVW�M�j���E �$���E�$���E�$�EP�MQ�M��ۂ��_^[��]�  ������������������������������U���DSVW�M��E�� ��E��@    �E��@    �E��@    �E�_^[��]��������������������U���DSVW�M��M��l����E��t�E�P�������E�_^[��]� ����������������������������U���DSVW�M��E�� ��E��x u�E��HQ�TZ	�B4��у��E��@    �E��@    _^[��]���������������������������������U���DSVW�M��EP�M��QR�TZ	�H4�Qt�҃�_^[��]� ����������������U���HSVW�M��} tB�EP�M�����P�TZ	�Q0���   �Ѓ��E��EP�M�Q�TZ	�B0���   �у���EP�M��QR�TZ	�H0�Q|�҃�_^[��]� ����������������������������������������U���DSVW�M��E��HQ�TZ	�B4�H�у�_^[��]����������������������U���DSVW�M��E��HQ�TZ	�B4�H�у�_^[��]����������������������U���DSVW�M��E��HQ�TZ	�B4�H�у�_^[��]����������������������U���DSVW�M��E��HQ�TZ	�B4�H|�у�_^[��]����������������������U���DSVW�M��E��HQ�TZ	�B4���   �у�_^[��]�������������������U���DSVW�M��E$P�M Q�UR�EP���E�$���E�$�M��QR�TZ	�H4��  �҃�$_^[��]�  �������������������������������U���DSVW�M��EP�MQ�UR�EP�M��QR�TZ	�H4�Q�҃�_^[��]� ��������������������U���DSVW�M��EP�MQ�UR�EP�M��QR�TZ	�H4�Q�҃�_^[��]� ��������������������U���DSVW�M��M�n�����u�M�gt��P�M��}����6�M�N�����u�M踣��P�M������hP�� A	��P��y����_^[��]� �������������������������������������U���DSVW�M��E�P�TZ	���   �B�Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	���   �B@�Ѓ�_^[��]����������������������U���DSVW�M��EP�M��QR�TZ	�H4�Q �҃�_^[��]� ����������������U���DSVW�M��EP�M��QR�TZ	�H4�Q$�҃�_^[��]� ����������������U���DSVW�M��EP�MQ�UR�EP�M��QR�TZ	�H0���   �҃�_^[��]� �����������������U���DSVW�M��EP�M��QR�TZ	�H0���   �҃�_^[��]� �������������U���DSVW�M����E�$�EP�MQ�U��BP�TZ	�Q0���   �Ѓ�_^[��]� �������������������������������U���DSVW�M��EP�M��QR�TZ	�H4���   �҃�_^[��]� �������������U���DSVW�M��EP�MQ�UR�EP�MQ�U��BP�TZ	�Q4���   �Ѓ�_^[��]� ����������������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U��BP�TZ	�Q4���   �Ѓ�_^[��]� ����������������������������U���DSVW�M��EP�M��QR�TZ	�H4�Q(�҃�_^[��]� ����������������U���DSVW�M��EP�MQ�UR�E��HQ�TZ	�B4�H,�у�_^[��]� �����������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4�B0�Ѓ�_^[��]� ���������������������������U���DSVW�M��E��HQ�TZ	�B4�H4�у�_^[��]����������������������U���hSVW�M��E�    �E�    �E�P�M�Q�UR�E��H�r����M��t���P�M��я���E�P�M�Q�U�R�E�P�M�Q�U��J��s���} tC�} t=�E�;E�~'�M�M�9M�}�U�;U�~�E�E�9E�}	�E�   ��E�    �E��V�.�} t(�E�;E�~�M�M�9M�}	�E�   ��E�    �E��&�E�;E�~�M�M�9M�}	�E�   ��E�    �E�_^[��]� �������������������������������������������������������������������������U���DSVW�M��EP�M��QR�TZ	�H4�Q8�҃�_^[��]� ����������������U���DSVW�M��EP�M��QR�TZ	�H4�Q<�҃�_^[��]� ����������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4���   �Ѓ�_^[��]� ������������������������U���DSVW�M����E�$�E��HQ�TZ	�B4��  �у�_^[��]� �����������������������U���DSVW�M��E��HQ�TZ	�B4�H@�у�_^[��]����������������������U���DSVW�M��E��HQ�TZ	�B4��  �у�_^[��]�������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4�BD�Ѓ�_^[��]� ���������������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4�BH�Ѓ�_^[��]� ���������������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4�BL�Ѓ�_^[��]� ���������������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4�BP�Ѓ�_^[��]� ���������������������������U���DSVW�M��M螏������   �M荏����u,�M�k��P�M�}k��P�E��HQ�TZ	�B4�HP�у��O�M�T�����u,�M辚��P�M�Dk��P�E��HQ�TZ	�B4�HH�у��hP��A	��P��p�����   �M� �������   �M������u,�M��j��P�M�P���P�E��HQ�TZ	�B4�HL�у��O�M趎����u,�M� ���P�M����P�E��HQ�TZ	�B4�HD�у��hP��A	��P�1p�����hP��A	��P�p����_^[��]� ��������������������������������������������������������������������������������������������U���DSVW�M��EP�MQ�UR�EP�M��QR�TZ	�H4��  �҃�_^[��]� �����������������U���DSVW�M��E,P�M(Q�U$R�E P�MQ�UR�EP�MQ�UR�EP�M��QR�TZ	�H4�QT�҃�,_^[��]�( ����������������������������U���DSVW�M��EP�MQ�UR�EP�M��QR�TZ	�H4�QX�҃�_^[��]� ��������������������U���DSVW�M��E��HQ�TZ	�B4�H`�у�_^[��]����������������������U���DSVW�M��E��HQ�TZ	�B4�Hd�у�_^[��]����������������������U���DSVW�M��EP�MQ�UR�EP�M��QR�TZ	�H4��   �҃�_^[��]� �����������������U���DSVW�M��EP�MQ�UR�EP�MQ�UR�E��HQ�TZ	�B4�H\�у�_^[��]� ���������������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4�Bh�Ѓ�_^[��]� ���������������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4��  �Ѓ�_^[��]� ������������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4��  �Ѓ�_^[��]� ������������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4�Bp�Ѓ�_^[��]� ���������������������������U���pSVW�M��E��x tp�} t(�M�����P�E��H�Ӂ��P�TZ	�Q0�Bl�Ѓ��B�M�����P�M��O���hARDb�M���t��P�E�P�M�Q�U��J�/q���M��ː���M��8l��_^[��]� ��������������������������������������������������U���DSVW�M��EP�M��QR�TZ	�H4�Ql�҃��   _^[��]� ���������������������������U���DSVW�M��EP���E�$���E�$�MQ�U��BP�TZ	�Q4���   �Ѓ�_^[��]� ����������������������U���DSVW�M��EP�MQ�UR�E��HQ�TZ	�B4���   �у�_^[��]� ��������������������U���DSVW�M��E��HQ�TZ	�B4���   �у�_^[��]�������������������U���DSVW�M��E��HQ�TZ	�B4��  �у�_^[��]�������������������U���DSVW�M��   _^[��]���������U���DSVW�M��   _^[��]���������U���DSVW�M�h�  �M��s���EP�MQ�UR�EP�M��u���2�_^[��]� ��������������������U���DSVW�M��EP�MQ�UR�EP�M���M��B��_^[��]� ��������������U���DSVW�M��   _^[��]� ������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�_^[��]� �����������U���DSVW�M�3�_^[��]� ���������U���DSVW�M�_^[��]� �����������U���DSVW�M��EP�MQ�UR�EP�M��QR�TZ	�H4�Qx�҃�_^[��]� ��������������������U���DSVW�M��EP�MQ�UR�E��H�b���_^[��]� ��������������������U���DSVW�M��} tj j�M�4���M��} tj j�M����M��EP�MQ�U��BP�TZ	�Q4�Bp�Ѓ�_^[��]� �����������������������������U���hSVW�M��E�    �M�o���E��}�INIbT�}�INIb��   �}�SACb,�}�SACb��   �}�$'  ��  �}�MicM��  ��  �}�ARDb��   �  �}�NIVb(�}�NIVbtJ�}�NPIb�:  �}�ISIb��   �~  �}�cnys�H  �l  �E���M��B���E�   �S  �E���M��B���E�   �:  �E�    �E�    �E�P�M�Q�U���M��P�҅�t �E�P�M�Q�U��BP�TZ	�Q4�B�Ѓ��E�   ��   �M��y��P�M��&q��P�E���M��B���E�   �   j j�M�X}���E�j j�M�I}���E�j j�M�:}���E�j j�M�+}���E܋EP�M�Q�U�R�E�P�M�Q�U���M��P���E�   �V�EP�M���M��B���F�EP�M���M��B$���E�   �)j hIicM�M��|���E��EP�M�Q�U���M��P ����E�_^[��]� ����������������������������������������������������������������������������������������������������������������������������������������������������������U���DSVW�M�h����h����h�����EP�MQh����h����h����h�����UR�M��c��_^[��]� ��������������������U���XSVW�M�hYALf�M��m��P�M���p���M��d��_^[��]����������������U���DSVW�M��M��^���E�� ���E��@   �E�_^[��]����������������U���DSVW�M��M��ˁ���E��t�E�P�i�����E�_^[��]� ����������������������������U���DSVW�M��E�� ���M��h|��_^[��]�������������U���HSVW�M��M�kk���E��}�cksat6�}�ckhct�G�E��@   �M��}����t�E��@    �   �03��,�E��x t�E���M��B���3���EP�MQ�M��p��_^[��]� �������������������������������������U���@SVW�EP�MQ�UR�EP�MQ�UR�TZ	�H���  �҃�_^[��]����������������������U���@SVW�EP�TZ	�Q0���   �Ѓ�_^[��]�������������������������U���PSVW�EP�MQ�U�R�TZ	�H0���   �҃�P�M覆���M���`���E_^[��]������������������������������U���|SVW�M�舂���E�    �	�E���E�   ����   j �E�k�
P�M��x���E�j �E�k�
��P�M�x���E�}� u�S�}� ~#j hе�M��}����E�P�M��m����M��9`���E�P�M�Q�U�R�[x����P�M��H����M��`���d����E�P�M赅���M���_���E_^[��]�������������������������������������������������������������U���DSVW�M�j�j��EP�M��o���P�M���y���E�_^[��]� ���������������U���@SVW�EP�MQ�TZ	�B0���   �у�_^[��]���������������������U���@SVW�EP�MQ�UR�EP�MQ�UR�TZ	�H0���   �҃�_^[��]����������������������U���@SVW�EP�TZ	�Q0���   �Ѓ�_^[��]�������������������������U���@SVWj0j 萄����P�EP�^����_^[��]������������������������U���@SVW�EE_^[��]�����������U���@SVWj0j �0�����P�EP�U\����P�'^����_^[��]���������������U���PSVWj0j �������P�EP�MQ�U�R�k����P��]�����M���]��_^[��]�������������������������������U���PSVWj0j 萃����P�EP�MQ�UR�E�P�h����P�{]�����M��f]��_^[��]���������������������������U���@SVWj j�0�����P�EP�0]����3Ƀ�����_^[��]��������������U���@SVWj j�������P�EP�[����P��\����3Ƀ�����_^[��]���������������������U���TSVWj j蠂����P�EP�MQ�U�R�bj����P�\����3Ƀ����M��M��o\���E�_^[��]���������������������������������U���TSVWj j�0�����P�EP�MQ�UR�E�P�7g����P�\����3Ƀ����M��M���[���E�_^[��]�����������������������������U���@SVW�EP�MQj �TZ	�B���   �у�_^[��]�������������������U���@SVW�EP�MQ�URj �TZ	�H���   �҃�_^[��]����������������U���DSVW�M��EP�MQ�UR�E��HQ�TZ	�B4�H,�у�_^[��]� �����������������������U���DSVW�M��EP�MQ�U��BP�TZ	�Q4�B0�Ѓ�_^[��]� ���������������������������U���DSVW�M��E��HQ�TZ	�B4�H4�у�_^[��]����������������������U���LSVW�M��M�x\��� �E��M�d���E�}� t�E�   �E�P�M�Q�UR�M��g��_^[��]� ����������������������������������U���DSVW�M��E P�MQ�M�gc��P�UR�EP�MQ�M��x���R�EP�M��|��_^[��]� �����������������������U���DSVW�M��M�w��P�E<P���E4�$���E,�$�M(Q���E �$���E�$���E�$�M�f����� �$�UR�M���e��_^[��]�8 ���������������������������������U���DSVW�M��M�w��P���E �$���E�$���E�$�M�9f����� �$�EP�M��g��_^[��]�  ���������������������������U���DSVW�M��M�v��P���E �$���E�$���E�$�M��e����� �$�EP�M��{��_^[��]�  ���������������������������U���DSVW�M��M�0v��P���E �$���E�$���E�$�M�Ye����� �$�EP�M��jh��_^[��]�  ���������������������������U���DSVW�M��M�)]��P�EP�MQ�UR�M��e��P�EP�MQ�M��'a��_^[��]� �����������������������������U���DSVW�M��EP�M��n��P�M�6e��P�MQ�M���m��_^[��]� �������������������������U���DSVW�M��E P���E�$���E�$�M�+g��P�MQ�M��)\��_^[��]� ����������������U���`SVW�M��E�P�M�Q�UR�M�胂���E�P�M�Q�U�R�E�P�MQ�M��V���} tC�} t=�E�;E�~'�M�M�9M�}�U�;U�~�E�E�9E�}	�E�   ��E�    �E��V�.�} t(�E�;E�~�M�M�9M�}	�E�   ��E�    �E��&�E�;E�~�M�M�9M�}	�E�   ��E�    �E�_^[��]� ��������������������������������������������������������������U���LSVW�M��E�E��}� u	�E����E�j hdiuM�M�m���E�}� u�   �G�E��M�;u3��9j hIicM�M�m��9E�uj h1icM�M�i����t3���E��M��   _^[��]� ������������������������������������������������U���DSVW�M��EP�MQ�TZ	�B�M����   ��_^[��]� ���������������U���XSVWhfnic�M�1g���E��}� tj
�M�誀����t�Vhfnic�E�P�M�X��P�M�_���M��U���M�f]�����t�M�Y]����uhfnic�M�O`���EPj
�M�L���_^[��]�������������������������������������U���DSVW�M��EP�TZ	�Q�M��B$��_^[��]� ����������������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���XSVW�M��EP�M�Q�TZ	�B�M��PP��P�M�=l���M��T���E_^[��]� ������������������������������U���DSVW�M��EP�TZ	�Q�M��BT��_^[��]� ����������������������U���DSVW�M��EP�MQ�UR�EP�M��^i��P�TZ	�Q0���   �Ѓ�_^[��]� ������������������������������U���DSVW�M��M�)l��Pj j j �EP�MQj �M�wd��Pj=�U��BP�TZ	�Q0���   �Ѓ�(_^[��]� ����������������������������U���DSVW�M��M�k��P�EPj j j��MQj �M�d��Pj=�U��BP�TZ	�Q0���   �Ѓ�(_^[��]� ����������������������������U���DSVW�M�j j j j j j j j j6�M��h��P�TZ	�H0���   �҃�(_^[��]��������������������������������U���HSVW�M�j �EP�M��f���E��E�P�M���N��_^[��]� ��������������U���HSVW�M�j �EP�M�i���E��E�P�M��m��_^[��]� ��������������U���LSVW�M������$�EP�M�qe���]���E��$�M��n��_^[��]� �������������������U���   SVW�M��M���n����t�����n��P�EP�M�Q�M�M����U�H�M�P�U�H�M��P�U�@�E����ċM��U�P�M�H�U��P�M�H�U��P�M��L��_^[��]� �������������������������������������������������U���tSVW�M��M��kp���M��cp��P�EP�M�Q�M�q����U�H�M��P�U�@�E����ċM��U��P�M�H�U��P�M���h��_^[��]� �������������������������������U���xSVW�M��M���p���M���p��P�EP�M�Q�M�)r��P�M���R���M���N���M���N�����̍E�P�st���M��k���M��N��_^[��]� �����������������������������������U���PSVW�M��E;Eu&j htsem�M�f����uj hrdem�M�f����t3��<�E�    �EP�M��i���M�Q�U�R�M�S����u3���E�P�M���K���   _^[��]� ���������������������������������������������U���PSVW�M��E;Eu&j htsem�M��e����uj hrdem�M��e����t3��<�E�    �EP�M���h���M�Q�U�R�M�Fv����u3���E�P�M��Rj���   _^[��]� ���������������������������������������������U���TSVW�M��E;Eu&j htsem�M�?e����uj hrdem�M�,e����t3��?���]�EP�M��$h���M�Q�U�R�M�by����u3�����E��$�M��j���   _^[��]� ������������������������������������������U���tSVW�M��E;Et�E;Et�E;Et3��   j htsem�M�xd����uj hrdem�M�ed����t3��   �����$�M��{[���EP�M��Og���MQ�M��Cg���UR�M��7g���E�P�M�Q�U�R�E�P�M�w����u3��5���ċM��U�P�M�H�U��P�M�H�U��P�M��=H���   _^[��]� ����������������������������������������������������������������������U���\SVW�M��E;Eu&j htsem�M�_c����uj hrdem�M�Lc����t3��Y�M���k���EP�M��Af���M�Q�UR�E�P�M��o����u3��)���ċM��U��P�M�H�U��P�M��:d���   _^[��]� ������������������������������������������������U���hSVW�M��E;Eu&j htsem�M�b����uj hrdem�M�|b����t3��d�M��l���EP�M��qe���M�Q�U�R�M�jM����u�E�    �M�� J���E��(���̍E�P�o���M��<f���E�   �M���I���E�_^[��]� �����������������������������������������������������U���DSVW�M��M���l���E�� ܵ�E��M�Hj hmyal�M�a���M��A�E��xt�E��xt
�E��@    j
hhfed�M�la���M��A�E�_^[��]� ����������������������������������������U���DSVW�M��M��*U���E��t�E�P�O�����E�_^[��]� ����������������������������U���DSVW�M��M��g��_^[��]����������������������U���HSVW�M��M�{Q���E��}�ytsdt��M��r���E���M��B�и   ��EP�MQ�M��i��_^[��]� �������������������������U���DSVW�M�3�_^[��]������������U���DSVW�M�3�_^[��]������������U���DSVW�M�_^[��]��������������U���DSVW�M�3�_^[��]������������U���DSVW�M�3�_^[��]������������U���DSVW�M�3�_^[��]������������U���DSVW�M�3�_^[��]� ���������U���\SVW�M��M��IF���E�P�M��W���M���E���E_^[��]� ����������������������������U���DSVW�M��M����l��_^[��]�������������������U���DSVW�M��E��M���E��P�M����*b���E�_^[��]� ����������������������������U���DSVW�M��E���M��BD�Ѕ�t!�E��H;Mt�E��M�H�E���M��BH��_^[��]� �������������������������U���DSVW�M��E��@_^[��]��������U���DSVW�M��E��x u3���E��H��������_^[��]����������������U���DSVW�M�_^[��]��������������U���DSVW�M��D�_^[��]���������U���DSVW�M������$�E��H�\���E�P�M��Q�E��H��B$��j j h����mk����_^[��]�����������������������������������U���DSVW�M��E��E�X(_^[��]� ������������������U���   SVW�M���T���P�M���M��B(��P�M���j����T����~D��j j j ��d����Af��Pj jj?j �M���A����d����QD��j ��x����f��Pj j(�`U����Pjh�  �M��Le���������w�����x����D����w�����t3��   j j j �M���e��Pj j j8j �M��^A���M���C��j�M��:I���M��{A��Pj��T����Ph,  ��T����Pj;�M��te��Ph	��h�  �M��"@���M��C���M���D���M��2E���M��*E��j�M���O���E��M��H$j�h`�����   _^[��]������������������������������������������������������������������������������������������������U���@SVWj �EP��H����_^[��]�������������������U���@SVW�E��E_^[��]��������U���\SVW�M�j�M����Oe���E��@4    �E��@8    �E��@<    �E����X(h�   �M��U��j hX��M��jg��h�  �M��{]��j j �E�P�M�Q�M���X���M��B��j j�M����HV��_^[��]���������������������������������������U���DSVW�M��E���_^[��]��������U���HSVW�M��E�    �   ����   �E��x4 t8hP��DA	��P�UB����j
�_�����M����nH����t3��   뿋M���0�w^���E��x4 ur�E��M�H8�E��M�H4�M���0�J���E��x4 tj
�;_�����M����H����t3��X�؋M���0�^���E��H<�M��E��@<    �M���0�I���(�!hP��DA	��$P�A�����M���0�I�������E�_^[��]� �����������������������������������������������������������������������U���DSVW�M��TZ	�PP�M��Bh��_^[��]��������������U���DSVW�M��TZ	�PP�M��Bl��_^[��]��������������U���DSVW�M��E��HQ�TZ	�BP�H�у�_^[��]����������������������U���   SVW�M�j h\���X�����d��h�  �M���Z��j j ��X���P�M��A(�H��M��P��h���R��b����P��x���P�wk����P�M�Q�M��V����x����3?����h����(?����X����?��htats�M���H��jj�M��lO���E����@(�$j�M��=��h�  �M��/Z���E�P�M�Q�U�R�M��E���M��d���E��x4 tc�M���0��[���E��x4 t.�E��H8Q�U��B4�Ѓ��M��A<�E��@8    �E��@4    �hP��HA	��P�C?�����M���0�<G���M��?��_^[��]� ���������������������������������������������������������������������������������������������������U���PSVW�EP�M��c���EP�M���f���E�P�M�jc���M��=���E_^[��]������������������U���   SVW�M��M�F����x�����x���MicMt}��x���ckhctM��x���fnict��   j��|����G��P�M�H����|����>��jj�M�S���   �   �   �E���M��B�Ѕ�u3��   �   �   �wj hIicM�M�U����x�����x������t�Thtats�M��F��j j�M��M��h�  �M���W���E�P�M�Q�U�R�M���B���M��}b���M���=��j�M��f���EP�MQ�M���_��_^[��]� ������������������������������������������������������������������������������������������U���HSVW�M��E�E��}�t�(j�M����^��j��X����j �M��Ue���   ��EP�MQ�M��G��_^[��]� �������������������������������������U���DSVW�M�j�M����?^��j�zX����3�_^[��]���������������������U���TSVW�M��M�����8���E�� �����M���8��P�M����8���M���`���E�_^[��]���������������������������U���DSVW�M��E��     �E��@    �E�_^[��]������������������������U���DSVW�M�j �E�P�M��a���E�_^[��]� ����������U���DSVW�M��EP�M�Q�UR�TZ	���   �Q�҃�_^[��]� ����������������������������U���DSVW�M��E�3Ƀ8����_^[��]�����������������U���DSVW�M��E���_^[��]��������U���DSVW�M��E��8�u�E��     �E��M�H��E��8 u�E��H;Mt	�E��    _^[��]� �������������������U���DSVW�M��E�3Ƀ8����_^[��]�����������������U���DSVW�M��E���_^[��]��������U���DSVW�M��E��8�u�E��     �EP�M����=���$�E��8 u�EP�M����sU����t	�E��    �M��8��_^[��]� �����������������������������U���DSVW�M��EP�M���7�������_^[��]� ���������U���DSVW�M��E�3Ƀ8����_^[��]�����������������U���DSVW�M��E���_^[��]��������U���DSVW�M��E��8�u�E��     �E��M�H��E��8 u�E��H;Mt	�E��    _^[��]� �������������������U���DSVW�M��E�3Ƀ8����_^[��]�����������������U���DSVW�M��E���_^[��]��������U���DSVW�M��E��8�u�E��     �E��E�X�#�E��8 u�E��@�E������D{	�E��    _^[��]� ����������������������������U���DSVW�M��E���_^[��]��������U���DSVW�M��E��8�u4�E��     �E����M��U�P�M�H�U�P�M�H�U�P�(�E��8 u �EP�M���Q�o3������t	�E��    _^[��]� ���������������������������������������U���DSVW�E�M� �������Dz3�U�E�B�@������Dz�M�U�A�B������Dz	�E�    ��E�   �E�_^[��]���������������������������������U���DSVW�M��E�3Ƀ8����_^[��]�����������������U���DSVW�M��E���_^[��]��������U���DSVW�M��E��8�u(�E��     �E����M��U�P�M�H�U�P�(�E��8 u �EP�M���Q��/������t	�E��    _^[��]� �����������������������������������U���LSVW�E�M� �������Dz�E�M�@�A������Dz3��T�E�M� �I���$�ca�����U�E��H���$�]��Ga�����E�������D{	�E�   ��E�    �E�_^[��]�������������������������������������������������U���`SVW�M�j h�  �M��R���} u�   �kj h�  �M��KE���E��}� u3��O�M��1���EPh�  �M��0D�����E�$h�  �M��E2��j �E�P�M��&C���E�   �M���4���E�_^[��]� ����������������������������������������������������U���DSVW�M��EP�MQ�U�R�TZ	�H@�Q(�҃�_^[��]� ���������������U���DSVW�M����E�$�E�P�TZ	�QH�B�Ѓ�_^[��]� �������������U���DSVW�M��EP�M�Q�TZ	�BH���   �у�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�BH���  �у�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�BH���  �у�_^[��]� ���������������U���DSVW�M��EP�MQ�U�R�TZ	�HH��  �҃�_^[��]� ����������������������������U���DSVW�M��EP�MQ�U�R�TZ	�HH��  �҃�_^[��]� ����������������������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�BH���  �у�_^[��]� ���������������U���DSVW�M�j �E�P�TZ	�QH���   �Ѓ�_^[��]��������������������U���DSVW�M��EPj �M�Q�TZ	�BH���   �у�_^[��]� �������������U���DSVW�M�j�E�P�TZ	�QH���   �Ѓ�_^[��]��������������������U���DSVW�M��EPj�M�Q�TZ	�BH���   �у�_^[��]� �������������U���DSVW�M�j�E�P�TZ	�QH���   �Ѓ������_^[��]��������������U���DSVW�M��EPj�M�Q�TZ	�BH���   �у�_^[��]� �������������U���DSVW�M��EP�MQ�U�R�TZ	�HH���   �҃�_^[��]� ����������������������������U���DSVW�M��EP�MQ�U�R�TZ	�HH���   �҃�_^[��]� ����������������������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�HH���  �҃�_^[��]� ����������������U���HSVW�M��EP��U�����E��}� t�EP�M�Q�M��-���E�_^[��]� �������������������U���HSVW�M��EP�MQ�RX�����E��}� t�EP�M�Q�M��k-���E�_^[��]� �������������������������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�BH���   �у�_^[��]� ���������������U���DSVW�M��EP�MQ�U�R�TZ	�HH���  �҃�_^[��]� ����������������������������U���DSVW�M��EP�M�Q�TZ	�BH���   �у�_^[��]� ���������������U���DSVW�M��EP�MQ�U�R�TZ	�HH��8  �҃�_^[��]� ����������������������������U���DSVW�M��EP�MQ�U�R�TZ	�HH��   �҃�_^[��]� ����������������������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH��  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH��  �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�U�R�TZ	�HH��  �҃�_^[��]� ����������������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QH��   �Ѓ�_^[��]� �����������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�BH��|  �у�_^[��]� �������������������U���DSVW�M��EP�M�Q�TZ	�BH��  �у�_^[��]� ���������������U���DSVW�M��E�P�TZ	�QH��T  �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�U�R�TZ	�HH��  �҃�_^[��]� ����������������������������U���DSVW�M��EP�M�Q�TZ	�BH��8  �у�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�BH��<  �у�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QH��@  �Ѓ�_^[��]� �����������������������U���DSVW�M��EP�M�Q�TZ	�BH���  �у�_^[��]� ���������������U���DSVW�M��E�P�TZ	�QH��L  �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�BH��H  �у�_^[��]� ���������������U���HSVW�M�j h�  �M��4�����0?���E��M���-�����}�u�E���3�_^[��]�������������������������U���DSVW�M��E�P�TZ	�Q@�B,�Ѓ�_^[��]�������������������������U���DSVW�M�h�  �M��$��_^[��]�����������������U���DSVW�M��EP�M�Q�TZ	�BH���   �у�_^[��]� ���������������U���DSVW�M�j h�  �M��C,�����;��_^[��]������������������������U���\SVW�M��EP�MQ���E�$�U�R�E�P�TZ	�QH��  �Ѓ��M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[��]� ��������������������������������������U���\SVW�M��EP�MQ���E�$�U�R�E�P�TZ	�QH��  �Ѓ��M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[��]� ��������������������������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QH��   �Ѓ�_^[��]� �����������������������U���@SVW�TZ	�HH��  ��_^[��]�����������������U���@SVW�EP�TZ	�QH��  �Ѓ�_^[��]�������������������������U���DSVW�M����E�$�E�P�TZ	�QH��$  �Ѓ�_^[��]� ��������������������������U���DSVW�M��E�P�TZ	�QH��(  �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�U�R�TZ	�HH��,  �҃�_^[��]� ����������������������������U���DSVW�M��EP���E�$�MQ�U�R�TZ	�HH��0  �҃�_^[��]� �������������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH��4  �Ѓ�_^[��]����������������������U���DSVW�M��E��     �E�_^[��]������������������U���DSVW�M�j�E��Q�TZ	�BH��|  �у�_^[��]������������������U���DSVW�M��EP�TZ	�QH��x  �Ѓ��M���E�3Ƀ8 ����_^[��]� �����������������U���DSVW�M�j �E��Q�TZ	�BH��|  �у�_^[��]������������������U���DSVW�M��E�P�TZ	�QH��P  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH��T  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH��X  �Ѓ�_^[��]����������������������U���\SVW�M��E�P�M�Q�TZ	�BH��\  �у��U��
�H�J�H�J�H�J�H�J�@�B�E_^[��]� �����������������������U���DSVW�M��E�P�TZ	�QH��`  �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�BH��d  �у�_^[��]� ���������������U���DSVW�M����E�$�E�P�TZ	�QH��h  �Ѓ�_^[��]� ��������������������������U���DSVW�M����E�$�E�P�TZ	�QH��t  �Ѓ�_^[��]� ��������������������������U���DSVW�M����E�$�E�P�TZ	�QH��l  �Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�M�Q�TZ	�BH��p  �у�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�BH���  �у�_^[��]� �������������������U���DSVW�M��EP�MQ�UR�EP�MQ�UR�E�P�TZ	�QH���  �Ѓ�_^[��]� ���������������������������U���@SVW�E P�MQ���E�$�UR�EP�MQ�TZ	�BH���   �у�_^[��]��������������������������������U���@SVW�EP���E�$�MQ�UR�EP�TZ	�QH���   �Ѓ�_^[��]��������������������U���@SVW�E�M�����*���E�EP�MQ�UR��C����_^[��]�������������������������U���@SVW�E;E}�E��E;E~�E��E_^[��]��������������������U����   SVW�M�1#���E��E�    �M�2���E��E�    �E�    �E�    �E�    �}� u
�   �H  �M�>��=�  �K	  j h:  �M�68���E؋M�)&���E��E�    �M�<���E��M�����E��M�5���E��E�    �	�E���E�E�;E���   �}� taj��E�P�M���=���EЃ}��tJ�M�k�M��_:��9E�t빋M�k�M������E��E�;E�~�E��EċM�k�M��m ��E��E��0�E����M����U��u��D;Du�E����E��	�E����E��O����}� tj �EP�M��(#����u
��  ��  �}� tn�M��?����tb�M���#��;E�uUhض�LA	��%P�M�k�Q�TZ	�B���  �у��E�}� u
�  �  �E�P�M�Q�M��)?��P�����hض�LA	��)P�M�k�Q�TZ	�B���  �у��E�}� u
�C  �>  �E�P�M�Q�U�R�\�����}� ~?hض�LA	��.P�M�����Q�TZ	�B���   �у��E܃}� u
��
  ��
  j��E�P�M�/����u
��
  ��
  �}� tj�EP�M���!����u
�
  �
  �}� t�M��d����<����
ǅ<���    ��<����E��M�0/���E��E�    �E�    �	�E���E�E�;E��m  �}� ��  j��E�P�M��;���EЃ}����  �M�k�M���7��9E�t뱋M�k�M��&���E��E�    �E�    �E�    �	�Ẽ��E̋M�k�M���5��9E��  �E�P�M�k�M��g6����u�ȋE�P�M�k�M������E��E����MȋU܋u�����Mȃ��MȋE����MȋU܉��Eȃ��EȋE����MȋU܋u��D���Mȃ��MȋE���   �UȋE܉��Mȃ��MȋE����MȋU܋u��D���Mȃ��MȋE���   �UȋE܉��Mȃ��MȋE����MȋU܋u��D���Mȃ��MȋE���   �UȋE܉��Mȃ��M�������EȉE��}� �
  �E��+���P�E�P�M��R���E�    �E�;E�|6hĶ�LA	��ZPhضh����3����hض�LA	��ZP������E�;E�|
�<  �7  �EȋM܋��U��}� t4�E�k�E�M�k�M����P�Q�P�Q�P�Q�P�Q�@�A�E�k�E�M�k�M���P�Q�P�Q�P�Q�P�Q�@�A�E�;E���   �EȋM܋�;U���   �EȋM܋D��������E��EȋM܋T����U��E���<�����<���wR��<����$����E����M��U���4�E����M��U��T�"�E����M��U��T��E����M��U��T�Eȃ��E��J����E����E��E����E��E�;E��b����E�;E�t6h���LA	��wPhضh���@2����hض�LA	��wP�x�����E�;E�t
�  �  �  �E����M����U��u��D3�;D�U��}� �  �E����M��k�U�E�k�E��
��J�H�J�H�J�H�J�H�R�P�E����M��Tk�U�E���k�E��
��J�H�J�H�J�H�J�H�R�P�E����M��Tk�U�E���k�E��
��J�H�J�H�J�H�J�H�R�P�}� tA�E����M��Tk�U�E���k�E��
��J�H�J�H�J�H�J�H�R�P�E����M��k�U�E�k�E�
��J�H�J�H�J�H�J�H�R�P�E����M��U���E����E��E����M��Tk�U�E�k�E�
��J�H�J�H�J�H�J�H�R�P�E����M��U��T�E����E��E����M��Tk�U�E�k�E�
��J�H�J�H�J�H�J�H�R�P�E����M��U��T�E����E��}� tY�E����M��Tk�U�E�k�E�
��J�H�J�H�J�H�J�H�R�P�E����M��U��T�E����E���E����M����U��u��D�D
�~����E�P��$�����E�P��$�����  �M�F5��=  ��  �M����E��M�x?���E��E�    �	�E���E�E�;E�}D�E�M��<� u��E�M��|� t�E�M����E��P�M���E�M����E��LP��M��hض�LA	�   P�M�k�Q�TZ	�B���  �у��E�}� u3��(  �E�P�M�Q�U�R� ����hض�LA	�   P�M���Q�TZ	�B���  �у��E��}� u3���  �E�P�M�Q�U�R��8�����E�+���P�E�P�M�Z����u�E�P�#�����E�P�#����3��  �M�'���E�M�3���E��E�    �E�    �E�    �	�E���E�E�;E���  �E�M��<� u���E�    �	�E����E��E����M�U�;���   �E���;E�}�E��M��T;U�|hض�LA	�   P������   �E�E�k�E�M�k�M���P�Q�P�Q�P�Q�P�Q�@�A�M����M��E��M��Tk�U�E�k�E�
��J�H�J�H�J�H�J�H�R�P�E����E��"����E�M��|� ��   �E���;E�}�E�E�;E�|hض�LA	�   P������   �E�E�k�E�M�k�M���P�Q�P�Q�P�Q�P�Q�@�A�M����M��E�k�E�M�k�M���P�Q�P�Q�P�Q�P�Q�@�A�M����M��E�M��U���U��!����E�    �	�E���E�E�+���9E�}�E�M��D�    �E�M���   �͍E�P�)!�����E�P�!�����   �&�E�P�
!�����E�P�� �����E�P�� ����3�_^[��]���0�B�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���DSVW�M��TZ	���   �M��B��_^[��]�����������U���DSVW�M��EP�MQ�U�R�TZ	�HH���   �҃�_^[��]� ����������������������������U���DSVW�M�j h�  �M����_^[��]���������������U���DSVW�M��EP�MQ�U�R�TZ	�HH���   �҃�_^[��]� ����������������������������U���DSVW�M�j h(  �M����_^[��]���������������U���DSVW�M�h(  �M����_^[��]�����������������U���DSVW�M�j h�  �M��4��_^[��]���������������U���DSVW�M�h�  �M��H��_^[��]�����������������U���DSVW�M��E��@_^[��]��������U���DSVW�M��E���U�����_^[��]� �����������U���DSVW�M��E�� %�����_^[��]�����������������U���DSVW�M��E���U���/��_^[��]� �����������U���DSVW�M��E�� %   ������_^[��]�������������U���HSVW�M��E��x ~�M��	�����E���E������E�_^[��]����������������������������U���TSVW�M��E�    �E�    �E�    �E�8 u'�MQ�M��x����uj�M��m����u	�E�    ��E�   �U�E���E�8 uc�M������} u�EP�MQ�UR�EP�MQ�M��E&���7�E�E���M���3���E�}� t�EP�MQ�UR�E�P�MQ�M��&���ыE�8 u�M��Q����t	�E�    ��E�   �M�U���E�8 u�M��$���EP�M��~%���   �M��G���} u�EPj �MQ�UR�EP�M��%���E��uh  �G*�����E��}� u3��^�M���P�M��,���E�E���M���2���E�}� t1�EPj �MQ�U�R�EP�M��4%���E��}� t�E�P�M����뾋E�_^[��]� ���������������������������������������������������������������������������������������������������������������������������U���DSVW�M��EP�TZ	���   �M��BH��_^[��]� �������������������U���DSVW�M��TZ	���   �M��Bx��_^[��]�����������U���DSVW�M��EP�TZ	���   �M��B|��_^[��]� �������������������U���DSVW�M��TZ	���   �M��B(��_^[��]�����������U���DSVW�M��EP�M�Q�TZ	�BH���   �у�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�BH���   �у�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�BH���   �у�_^[��]� ���������������U���DSVW�M��E�P�MQ�UR�TZ	�HH���   �҃�_^[��]� ����������������������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�U�R�TZ	�HH���   �҃�_^[��]� ����������������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�HH���  �҃�_^[��]� ����������������U���DSVW�M��E�P�TZ	�QH��t  �Ѓ�_^[��]����������������������U���DSVW�M��E�� 4��E��@    �E�_^[��]������������������������U���DSVW�M��M��w���E��t�E�P�������E�_^[��]� ����������������������������U���DSVW�M��E�� 4��E��HQ�TZ	�Bl�H�у�_^[��]�����������������������������U���DSVW�M��E��HQ�TZ	�Bl�H�у��} u�   �4�EP�MQ�UR�EP�TZ	�Ql��Ѓ��M��A�E�3Ƀx ����_^[��]� ����������������������������������U���DSVW�M��E��x u3���E��HQ�TZ	�Bl�H�у�_^[��]�������������������������U���LSVW�M��E�P�M�Q�UR�EP�M������E�;Eu�E����E�;Eu�E�����_^[��]� ��������������������U���DSVW�M��EP�MQ�UR�EP�M��QR�TZ	�Hl�Q�҃�_^[��]� ��������������������U���@SVW�EP���E�$�MQ�UR�TZ	�HH���  �҃�_^[��]�������������������������U���@SVW�EP�MQ�UR�EP�TZ	�QH���  �Ѓ�_^[��]�����������������������������U���@SVW�E P�MQ�UR�EP�MQ�UR�EP�TZ	�QH���  �Ѓ�_^[��]�����������������U���@SVW�E0P���E(�$�M$Q�U R�EP�MQ�UR�EP�MQ�UR�TZ	�HH���  �҃�,_^[��]���������������������������������U���@SVW�EP�MQ�UR�TZ	�HH���  �҃�_^[��]������������������U���DSVW�M��EP���E�$�M�Q�TZ	�BH���  �у�_^[��]� ����������������������U���HSVW�M��E�    �}u�M�����E��$�} u�M��1���E���}u�M������E��}� u3���E�P�MQ�M��0��_^[��]� �����������������������������������U���dSVW�M��p���E��}� t�} u3���   �M��R���E�M�������E��}� u�E���   �E�    �	�E���E�M���9E���   �E�P�M�Q�U�R�E�P�M�+����u�ȋE�E��	�E���E�E�;E�_�E����u$�E������M������U�u�D;Du���E���P�M�0����M���T��U܃}��t�E�P�M������K����E�_^[��]� ������������������������������������������������������������������������U���DSVW�M�j h�  �M���"��_^[��]���������������U���DSVW�M��EP�MQ�U�R�TZ	�HH��p  �҃�_^[��]� ����������������������������U���DSVW�M��EP�M��QR�TZ	�Hl�Q�҃�_^[��]� ����������������U���TSVW�M��M��M���E��}� u3��G  �E�    �}u�M������E��$�} u�M��i ���E���}u�M��0���E�}� u3���   �M������E�    �	�E����E��M����9E���   �E�P�M�P����E�}� u�ϋE�HQ�M�n�����t�E���P�M��$����E�HQ�M�L�����t�E���   Q�M�������E����M����U��u��D;Dt&�E�HQ�M�
�����t�E���   Q�M������E�HQ�M�������t�E���   Q�M����������   _^[��]� ������������������������������������������������������������������������������������������������������������U���DSVW�M��EP�M�Q�TZ	�B\�H,�у�_^[��]� ������������������U���@SVW�E P�MQ�UR�EP�MQ�UR�EP�TZ	�QH���   �Ѓ�_^[��]�����������������U���DSVW�M��E�P�TZ	�QH���   �Ѓ�_^[��]����������������������U���@SVW�EP�MQ�UR�EP�MQ�TZ	�BH���  �у�_^[��]�������������������������U���@SVW���E�$���E�$�����$�EP�M������$�
�����$�MQ�M����_^[��]������������������������������U���@SVW�E�]����Au�E��E�]����z�E��E_^[��]��������������������������U���   SVW��x������P�EP�M�Q�M�S������E�$���E�$���E��$�	�����$���E�$���E�$���E��$�	�����$���E�$���E�$���E��$�r	�����$�M����P�EP�M�]��_^[��]�����������������������������������������������������������U���@SVW�EP�TZ	�QH��Ѓ�_^[��]�������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVWh�  �TZ	�HH��҃�_^[��]�������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���DSVWh  ������E��}� u3��kj �EPh�  �M��� ����u�.�,j �EPh(  �M��� ����u��j j�M��q���E��$�}� t�E�P�TZ	�Q@�B�Ѓ��E�    3�_^[��]��������������������������������������������U���DSVW�M��EP�MQ�TZ	���   �M��P��_^[��]� ���������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���DSVWh�  �������E��}� u3��9�EP�MQ�M��B
����u"�}� t�E�P�TZ	�Q@�B�Ѓ��E�    �E�_^[��]������������������������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVW�EP�MQ�TZ	�BH�H�у�_^[��]������������������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���DSVW�M��EP�M�Q�TZ	�BH���  �у�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�BH���  �у�_^[��]� ���������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���@SVW�EP�MQ�TZ	�BH���  �у�_^[��]���������������������U���@SVW�E0P�M,Q�U(R�E$P�M Q���E�$���E�$�UR�EP�TZ	�QH��P  �Ѓ�,_^[��]�������������������������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�U�R�TZ	�HH���  �҃�_^[��]� ����������������������������U���DSVW�M��E�P�TZ	�QH��  �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QH���  �Ѓ�_^[��]� �����������������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QH���  �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�BH��  �у�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�BH��  �у�_^[��]� ���������������U���DSVW�M��E�_^[��]�����������U���DSVW�M�_^[��]��������������U���@SVW�TZ	�HH���  ��_^[��]�����������������U���@SVW�EP�TZ	�QH���  �Ѓ�_^[��]�������������������������U���DSVW�M��E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R�TZ	�HH���  �҃�0_^[��]�, ������������������������U���DSVW�M��E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�U�R�TZ	�HH���  �҃�0_^[��]�, ������������������������U���DSVW�M��E�P�TZ	�QH��,  �Ѓ�_^[��]����������������������U���DSVW�M��EP�M�Q�TZ	�BH��X  �у�_^[��]� ���������������U���DSVW�M��E�P�TZ	�QH��\  �Ѓ�_^[��]����������������������U���@SVW�EP�MQ�UR�EP�MQ�TZ	�BH��0  �у�_^[��]�������������������������U���@SVW�Ek�P�MQ�UR�����_^[��]����������U���DSVW�M��}~�EP�MQ�UR�M�����_^[��]� �����������������U���@SVW�E��P�MQ�UR� ����_^[��]����������U���LSVW�M��EP�MQ�f������tQhP�h}  hH�h@�hH��f�����P�������Ph   @j�M����P��������Z	��t��G�E�M���U�EP�M�������P�M�Q�UR�E�P�M�����EP�M�Q�UR�E�P�M�����_^[��]� ���������������������������������������������������������������U���@SVW�EE_^[��]�����������U���DSVW�EP�r�����;Ev�M�M���U�U��E�_^[��]���������������U���@SVW�E�M�3�;��_^[��]������������������U���HSVW�M��E�    ��E���E�}t�E����E���E�_^[��]� ����������������������U���LSVW�M��E+E���� ��   �} u�EP�MQ�UR�M������v�E���E�E��P�E+E���+����M��R�EP�MQ�M�������E��E�P�MQ�UR�EP�M�������E�EP�MQ�U�R�EP�M�����E�E�\���_^[��]� �������������������������������������������������������U���HSVW�M��} ~5�E   �E��E�P�MQ�UR�M�����EP�M�Q�UR�M��������E;Et�EP�MQ�UR�M�����_^[��]� ������������������������������������U���DSVW�M��EP�MQ��������t;�EP�MQ���������t�E�Y��EP�MQ���������t�E�>�E�9�4�EP�MQ��������t�E���EP�MQ��������t�E��E_^[��]� �����������������������������������������������������U���\�B	3ŉE�SVW�M��E+E���� ~�E+E��P�MQ�UR�M������   �E���E�E�E��E����E���E����E��M���M�E�;EtL�E�P�M�Q���������t8j�E�P�M�Q������j�E�P�M�Q������j�E�P�M�Q������뚋E���E�E�;E�t���_^[�M�3�������]� ���������������������������������������������������������������������U���P�B	3ŉE�SVW�M��E���E�   ����   �E���E�MQ�UR���������t��E���E�MQ�UR��������t��E;Er�E�Yj�EP�M�Q������j�EP�MQ������j�E�P�MQ�{������E;Eu�E�E��E;Eu�E�E�O���_^[�M�3�������]� �������������������������������������������������������������U���DSVW�M��	�E���E�E;Et�EP�MQ�M�������_^[��]� ����������������������U���l�B	3ŉE�SVW�M��}}�Z  �E�E�E�+������E�   ���9  �}�~�E���E��c�E���E�E�M�T���U�E�M���U�j�E�P�M�Q�1�����j�E�P�M�Q������j�E�P�M�Q�������}���   �E�E܋E܋M�T���U؋E���;E���   �E؉EԋE����E܋E܋M�T���U؋E�;E�})�E؃�P�M�Q��������t�E܃��E܋E؃��E؋E�P�M�Q��������t8j�E�P�M�Q�o�����j�E�P�M�Q�]�����j�E�P�M�Q�K��������S�������_^[�M�3������]� ������������������������������������������������������������������������������������������������������������������U���T�B	3ŉE�SVW�M��E��P�MQ��������t_j�EP�M�Q�y������E��E�j�E��P�MQ�^������E���E�E��P�M�Q�<�������u�j�E�P�MQ�,�����_^[�M�3������]� �������������������������������������������������U���HSVW�M��E�M��;t3���   �E�x uE�E�8 u=�E�x u4�E��x u�M��9 u�U��z u	�E�   ��E�    �E��   �I�E��x u@�E��8 u8�E��x u/�E�x u�M�9 u�U�z u	�E�   ��E�    �E��M�E�x t�E��x t�E�M��P;Qt3��)�E�x t�E��x t�E�M��P;Qt3���   _^[��]� ��������������������������������������������������������������������U���DSVW�M��EP�M�����������_^[��]� ������������������������U���HSVW�M��E�    �	�E����E��E�P�M������8 t��E�_^[��]����������������������U���LSVW�M��E�    �	�E����E��E�P�M�������8 t(�E�P�M����P�M�Q�M��������
����t�뾃} t�E�M���}� ~�E�P�M��s����8 u	�E�   ��E�    �E�_^[��]� ����������������������������������������U���DSVWj�P   ���E��}� t	�E��x u3���EP�MQ�UR�E��H�у�_^[��]��������������������������U���@SVWh\Z	�EPhD �����_^[��]�����������U���HSVW�M�j\�������E��}� t	�E��x\ u��E�P�M��Q\�҃��E�_^[��]������������������������������U���HSVW�M�j\�]������E��}� t	�E��x\ u��E�P�M��Q\�҃��EP�M��
���E�_^[��]� �������������������������������U���HSVW�M�j\��������E��}� t	�E��x\ u��E�P�M��Q\�҃��EP�M�������E�_^[��]� �������������������������������U���TSVW�M�j\�}������E��}� t	�E��x\ u�$�E�P�M��Q\�҃��EP�M��*���P�M��J����E�_^[��]� ����������������������U���DSVW�M��E��M��E��@    �E��@    �E�_^[��]� ����������������������������U���HSVW�M�j\�������E��}� t	�E��x\ u�'�E�P�M��Q\�҃��EP�M������EP�M��,����E�_^[��]� �����������������������������������U���HSVW�M�j\�=������E��}� t	�E��x\ u�3�E�P�M��Q\�҃��EP�M������EP�M������EP�M������E�_^[��]� ���������������������������������������U���HSVW�M�j`�������E��}� t	�E��x` u��E�P�M��Q`�҃�_^[��]�����������������U���HSVW�M�jd�]������E��}� t	�E��xd u��EP�M�Q�U��Bd�Ѓ�_^[��]� ��������������������������U���HSVW�M�jh��������E��}� t	�E��xh u��EP�M�Q�U��Bh�Ѓ�_^[��]� ��������������������������U���HSVW�M�jl�������E��}� t	�E��xl u��E�P�M��Ql�҃�_^[��]�����������������U���HSVW�M�h�   �J������E��}� t�E����    u3���EP�M�Q�U����   �Ѓ�_^[��]� �������������������������������U���HSVW�M�h�   ��������E��}� t�E����    u3���EP�M�Q�U����   �Ѓ�_^[��]� �������������������������������U���HSVW�M�jp�m������E��}� t	�E��xp u�`Z	��EP�M�Q�U��Bp�Ѓ�_^[��]� ���������������������U���PSVW�M�jt�������E��}� t	�E��xt uh`Z	�M�����E�+�EP�M�Q�U�R�E��Ht�у�P�M�'����M��&����E_^[��]� ����������������������������������U���HSVW�M�jx�}������E��}� t	�E��xx u�E���E�P�MQ�U��Bx�Ѓ��E�_^[��]� ��������������������U���HSVW�M�j|�������E��}� t	�E��x| u3���E�P�MQ�U��B|�Ѓ�_^[��]� ������������������������U���HSVW�M�j|�������E��}� t	�E��x| u�   ��E�P�MQ�U��B|�Ѓ������_^[��]� ������������������������������U���PSVW�M�h�   �J������E��}� t�E����    u�E��%�EP�M�Q�U�R�E����   �у��M��s����E�_^[��]� �������������������������������U���DSVW�M��E�_^[��]�����������U���DSVWj�������E��}� t	�E��x u3���E��H��_^[��]�������������������������U���DSVW�E�8 u�6j�V������E��}� t	�E��x u��EP�M��Q�҃��E�     _^[��]���������������������������������U���HSVW�M��} u3��7j��������E��}� t	�E��x u3���EP�MQ�U�R�E��H�у�_^[��]� ��������������������������U���HSVW�M�j�}������E��}� t	�E��x u3���EP�M�Q�U��B�Ѓ�_^[��]� ������������������������U���HSVW�M�j�������E��}� t	�E��x u3���EP�M�Q�U��B�Ѓ�_^[��]� ������������������������U���HSVW�M�j �������E��}� t	�E��x  u3���E�P�M��Q �҃�_^[��]�������������������������������U���HSVW�M�j$�]������E��}� t	�E��x$ u3���E�P�M��Q$�҃�_^[��]�������������������������������U���HSVW�M�j(��������E��}� t	�E��x( u3���EP�MQ�UR�E�P�M��Q(�҃�_^[��]� ��������������������������������U���HSVW�M�j,�������E��}� t	�E��x, u3���EP�MQ�U�R�E��H,�у�_^[��]� ��������������������U���HSVW�M�j(�-������E��}� t	�E��x0 u3���EP�MQ�UR�E�P�M��Q0�҃�_^[��]� ��������������������������������U���HSVW�M�j4�������E��}� t	�E��x4 u3���E�P�M��Q4�҃�_^[��]�������������������������������U���HSVW�M�j8�]������E��}� t	�E��x8 u3���EP�MQ�UR�EP�M�Q�U��B8�Ѓ�_^[��]� ����������������������������U���HSVW�M�j<��������E��}� t	�E��x< u��EP�M�Q�U��B<�Ѓ�_^[��]� ��������������������������U���HSVW�M�jD�������E��}� t	�E��xD u3���E�P�M��QD�҃�_^[��]�������������������������������U���HSVW�M�jH�-������E��}� u��EP�M�Q�U��BH�Ѓ�_^[��]� �������������������U���HSVW�M�jL��������E��}� u3���EP�M�Q�U��BL�Ѓ�_^[��]� �����������������U���HSVW�M�jP�������E��}� u3���EP�MQ�U�R�E��HP�у�_^[��]� �����������������������������U���HSVW�M�jT�-������E��}� u3���E�P�M��QT�҃�_^[��]������������������������U���HSVW�M�jX��������E��}� u��EP�M�Q�U��BX�Ѓ�_^[��]� �������������������U���HSVW�M�h�   �������E��}� u3��&�EP�MQ�UR�EP�MQ�U�R�E����   �у�_^[��]� ���������������������������U���HSVW�M�h�   �������E��}� u3���EP�MQ�UR�E�P�M����   �҃�_^[��]� �������������������U���HSVW�M�h�   �������E��}� u3���EP�M�Q�U����   �Ѓ�_^[��]� ���������������������������U���HSVW�M�h�   �Z������E��}� u3���EP�M�Q�U����   �Ѓ�_^[��]� ���������������������������U���HSVW�M�h�   ��������E��}� u3���EP�M�Q�U����   �Ѓ�_^[��]� ���������������������������U���HSVW�M�h�   �������E��}� u��EP�MQ�UR�E�P�M����   �҃�_^[��]� ���������������������U���TSVWh�   �=������E��}� u�M������E�*�EP�M�Q�U����   �Ѓ�P�M�����M�������E_^[��]������������������������������������U���LSVWh�   �������E��}� t�E����    u�EP�M������E�.�EP�MQ�U�R�E����   �у�P�M������M�������E_^[��]��������������������������������U���\SVW�M�h�   �*������E��}� t�E����    uj �M������P�M�"����E�*�EP�M�Q�U��M����   ��P�M�<����M��;����E_^[��]� ���������������������������������������U���HSVW�M�h�   �������E��}� t�E����    u3���EP�MQ�UR�E��M����   ��_^[��]� ���������������������������U���HSVW�M�h�   �������E��}� t�E����    u3���EP�U��M����   ��_^[��]� �������������������U���HSVW�M�h�   �������E��}� t�E����    u3���EP�U��M����   ��_^[��]� �������������������U���HSVW�M�h�   �Z������E��}� t�E����    u3���EP�U��M����   ��_^[��]� �������������������U���HSVW�M�h�   ��������E��}� t�E����    u3���E��M����   ��_^[��]��������������������������U���HSVW�M�h�   �������E��}� t�E����    u3���EP�MQ�UR�E��M����   ��_^[��]� ���������������������������U���HSVW�M�h�   �*������E��}� t�E����    u��EP�U��M����   ��_^[��]� ���������������������U���HSVW�M�h�   ��������E��}� t�E����    u3���EP�MQ�UR�E��M����   ��_^[��]� ���������������������������U���LSVW�M�h�   �Z������E��}� t�E����    u3���E��M����   �҉E�E�_^[��]��������������������U���DSVWj�`   ���E��}� t	�E��x u����'�E P�MQ�UR�EP�MQ�UR�EP�M��Q�҃�_^[��]�������������������������U���@SVWhpZ	�EPh�f ������_^[��]�����������U���PSVWj��������E��}� t	�E��x u�E������M�n����E��?�E8P�M4Q�U0R�E,P�M(Q���̍UR�����EP�M��Q�҃�4�E��M�-����E�_^[��]����������������������������������U���DSVWj� ������E��}� t	�E��x u3���EP�MQ�U��B�Ѓ�_^[��]������������������������������U���DSVWj��������E��}� t	�E��x u3���EP�M��Q�҃�_^[��]������������������U���DSVW�M��E�� ���E�_^[��]������������������U���DSVW�M��M��#����E��t�E�P�������E�_^[��]� ����������������������������U���DSVW�M��E�� ��_^[��]���������������������U���TSVW�M��E��E��}� t,�E��E��M��M��}� tj�U���M���҉E���E�    �E�    _^[��]�������������������������������U���DSVW�M��TZ	�P�M���  ��_^[��]�����������U���DSVW�M��TZ	�P�M���(  ��_^[��]�����������U���`SVW�M��E�P�TZ	�Q�M���   ��P�M�s����M������E_^[��]� �������������������������������U���DSVW�M��TZ	�P�M���$  ��_^[��]�����������U���@SVW�EP�MQ�TZ	�B��  �у�_^[��]���������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�TZ	�H��  ��_^[��]�����������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�TZ	�B��x  �у�_^[��]���������������������U���@SVW�EP�TZ	�Q��|  �Ѓ�_^[��]�������������������������U���@SVW�TZ	�H��d  ��_^[��]�����������������U���@SVW�EP�MQ�TZ	�B��p  �у�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B��t  �у�_^[��]���������������������U���HSVW�M��E�P�TZ	���   �BX�Ѓ��E��}� u3���EP�MQ�M��{���_^[��]� ����������������������U���DSVW�M��EP�MQ�U�R�TZ	�H|�Q�҃�_^[��]� ���������������U���HSVW�M��E�P�TZ	���   �BX�Ѓ��E��}� u3���EP�MQ�M�����_^[��]� ����������������������U���DSVW�M��EP�MQ�U�R�TZ	�H|�Q8�҃�_^[��]� ���������������U���DSVW�M��E��M�j j j �E��Q�TZ	�B�H�у��U��B�E�_^[��]� �����������������������������U���DSVW�M�j j j �E��Q�TZ	�B�H�у��U��B_^[��]���������������������������U���DSVW�M��E��x u3��0�E��HQ�UR�EP�M��R�TZ	�H�Q�҃��M��A�   _^[��]� ������������������������������U���DSVW�M�j j��TZ	�P�M��B�ЋE�_^[��]�����������������������U���DSVW�M�j �EP�TZ	�Q�M��B�ЋE�_^[��]� �����������������U���DSVW�M��EPj��TZ	�Q�M��B�ЋE�_^[��]� �����������������U���DSVW�M��M������_^[��]����������������������U���DSVW�M��TZ	�P�M��B��_^[��]��������������U���DSVW�M�j j �E�P�M�����E�_^[��]� ������������������������U���DSVW�M��EP�MQ�UR�TZ	�P�M����   ��_^[��]� ����������������������������U���DSVW�M��EP�M�Q�TZ	�B�H�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�B�H�у������_^[��]� ���������������������������U���HSVW�M��EP�M������E��M�����_^[��]� ��������������������U���DSVW�M��E�P�TZ	���   �BX�Ѓ�_^[��]����������������������U���DSVW�M��EP�TZ	�Q�M��Bt��_^[��]� ����������������������U���DSVW�M�h#  �EP�MQ�M��m���_^[��]� ����������������������U���DSVW�M��EP�MQ�UR�TZ	�P�M��Bl��_^[��]� ���������������U���DSVW�M�hF  �EP�MQ�M�����_^[��]� ����������������������U���HSVW�M��EP�M������E��EP�M�蔻��_^[��]� ����������������U���DSVW�M��EP�M�Q�TZ	���   �H`�у�_^[��]� ���������������U���DSVW�M��EP�TZ	�Q�M����   ��_^[��]� �������������������U���HSVW�M��EP�TZ	�Q�M����   �ЉE��}� u3���M������_^[��]� ������������������������������U���DSVW�M��EP�M�Q�TZ	�B8�HD�у�_^[��]� ������������������U���@SVW�TZ	�H8�Q<��_^[��]��������������������U���@SVW�E�Q�TZ	�B8�H@�у��E�     _^[��]�����������������U���@SVW�TZ	�H8���_^[��]���������������������U���@SVW�E�Q�TZ	�B8�H�у��E�     _^[��]�����������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q8�B�Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�MQ�U�R�TZ	�H8�Q�҃�_^[��]� ���������������U���DSVW�M��E�P�TZ	�Q8�B�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�B8�H �у�_^[��]� ������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�H8�Q$�҃�_^[��]� �������������������U���DSVW�M��EP�MQ�UR�EP�MQ�UR�E�P�TZ	�Q8�B�Ѓ�_^[��]� ������������������������������U���DSVW�M��EP�MQ�U�R�TZ	�H8�Q(�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q8�B,�Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q8�B�Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�H8�Q�҃�_^[��]� �������������������U���DSVW�M��EP�MQ�U�R�TZ	�H8�Q0�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Q8�B4�Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�M�Q�TZ	�B8�H8�у�_^[��]� ������������������U���@SVW�EP�MQ�UR�EP�TZ	�Q��x  �Ѓ�_^[��]�����������������������������U���@SVW�EP�MQ�TZ	�B��|  �у�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B���  �у�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B���  �у�_^[��]���������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q�B,�Ѓ�_^[��]������������U���@SVW�E P�MQ�UR�EP�MQ�UR�EP�TZ	�Q���  �Ѓ�_^[��]�����������������U���PSVW�M������E�P�TZ	�Q�B8�Ѓ��E�P�M�e����M�諴���E_^[��]�����������������������������U���@SVW�TZ	�H�Q<��_^[��]��������������������U���@SVW�EP�MQ�TZ	�B�H@�у�_^[��]������������������������U���@SVW�TZ	�H�QD��_^[��]��������������������U���@SVW�TZ	�H�QH��_^[��]��������������������U���@SVW�EP�MQ�UR�TZ	�H�QL�҃�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B�HP�у�_^[��]������������������������U���@SVW�EP�TZ	�Q��<  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q��,  �Ѓ�_^[��]�������������������������U���@SVW�E��PP�M��@Q�U��0R�E�� P�M��Q�UR�EP�TZ	�Q���   �Ѓ�_^[��]����������������������������������U���@SVW�TZ	�H���   ��_^[��]�����������������U���@SVW�TZ	�H���  ��_^[��]�����������������U���@SVW�EP�MQ�UR�EP�MQh�6  �TZ	�B���   �у�_^[��]��������������������U���@SVW�EP�TZ	�Q�B�Ѓ�_^[��]������������U���@SVW�EP�TZ	�Q��\  �Ѓ�_^[��]�������������������������U���`SVW�EPj hķ�M��9���P�M�Q�(������M�������E�P�TZ	�Q�B�Ѓ��M��װ��_^[��]����������������������������U���@SVW�EP�TZ	�Q�BT�Ѓ�_^[��]������������U���@SVW�EP�TZ	�Q�BX�Ѓ�_^[��]������������U���@SVW�EP�TZ	�Q�B\�Ѓ�_^[��]������������U���@SVW�TZ	�H�Q`��_^[��]��������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�TZ	�H�Qd��_^[��]��������������������U���@SVW�TZ	�H�Qh��_^[��]��������������������U���@SVW�EP�TZ	�Q�Bl�Ѓ�_^[��]������������U���@SVW�EP�TZ	�Q�Bp�Ѓ�_^[��]������������U���@SVW�EP�MQ�UR�TZ	�H�Qt�҃�_^[��]���������������������U���@SVW�EP�TZ	�Q��D  �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�UR�EP�TZ	�Q��  �Ѓ�_^[��]�����������������������������U���@SVW�EP�MQ�TZ	�B�Hx�у�_^[��]������������������������U���@SVW�EP�MQ�TZ	�B��@  �у�_^[��]���������������������U���\SVW�M��R����E�P�MQ�TZ	�B�H|�у��E�P�M�����M�贵���E_^[��]�������������������������U���@SVW�EP�MQ�TZ	�B���   �у�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B��h  �у�_^[��]���������������������U���@SVW�EP�MQ�UR�EP�TZ	�Q��d  �Ѓ�_^[��]�����������������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�TZ	�H���   ��_^[��]�����������������U���@SVW�EP�MQ�TZ	�B��l  �у�_^[��]���������������������U���@SVW�EP�TZ	�Q��   �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�UR�TZ	�H��  �҃�_^[��]������������������U���TSVW�M������E�P�TZ	�Q���   �Ѓ��E�P�M�����M��p����E_^[��]��������������������������U���@SVW�TZ	�H��`  ��_^[��]�����������������U���@SVW�EP�TZ	�Q��  �Ѓ�_^[��]�������������������������U���XSVW�EP�M�Q�TZ	�B���   �у��U��
�H�J�H�J�H�J�H�J�@�B�E_^[��]�����������������������������U���@SVW�EP�MQ�TZ	�B���  �у�_^[��]���������������������U���@SVW�EP���E�$���E�$�MQ�TZ	�B���   �у�_^[��]�������������������U���@SVW�EP�MQ�UR�TZ	�H���   �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���   �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���   �҃�_^[��]������������������U���@SVW�EP�MQ�TZ	�B���   �у�_^[��]���������������������U���@SVW�EP�MQ�TZ	�B���   �у�_^[��]���������������������U���@SVW�EP�TZ	�Q���   �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q���   �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q���   �Ѓ�_^[��]�������������������������U���PSVW�M��E�P�M�Q�U�R�E�P�TZ	�Q���   �Ѓ���u3���E�_^[��]�������������������������������U���PSVW�M��E�P�M�Q�U�R�E�P�TZ	�Q���   �Ѓ���u3���E�_^[��]�������������������������������U���PSVW�M��E�P�M�Q�U�R�E�P�TZ	�Q���   �Ѓ���u3���E�_^[��]�������������������������������U���@SVW�EP�TZ	�Q��8  �Ѓ�_^[��]�������������������������U���DSVW�M��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�λ��P�U�R�TZ	�H0���   �҃�(_^[��]�$ ���������������������������U���DSVW�M��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�M�"���P�U�R�TZ	�H0���   �҃�(_^[��]�$ ���������������������������U���DSVW�M��E��@_^[��]��������U���DSVW�M��E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�E�P�TZ	�Q0���   �Ѓ�(_^[��]�$ �������������������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�B0���   �у�_^[��]� �������������������U���DSVW�M��E�P�TZ	�Q0���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�U�R�TZ	�H0���   �҃�_^[��]� ����������������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�B0���   �у�_^[��]� �������������������U���DSVW�M��E�P�TZ	�Q0���   �Ѓ�_^[��]����������������������U���@SVW�TZ	�H0���   ��_^[��]�����������������U���@SVW�E�Q�TZ	�B0���   �у��E�     _^[��]��������������U���@SVW�EP�TZ	�Q��H  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q��T  �Ѓ�_^[��]�������������������������U���@SVW�TZ	�H��p  ��_^[��]�����������������U���@SVW�TZ	�H���  ��_^[��]�����������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�UR�EP�TZ	�Q���  �Ѓ�_^[��]�����������������������������U���@SVW�EP�MQ�UR�EP�MQ�TZ	�B���  �у�_^[��]�������������������������U���PSVW�EP�MQ�UR�E�P�TZ	�Q��X  �Ѓ�P�M�<����M��z����E_^[��]�������������������������U���dSVWj hLGOg�M�� ���PhicMC�E�P蠿�����M�蛠���M�萨����u�M�֜���M��
����E��M��o���P�M������M�������E_^[��]�������������������������������������������U���@SVW�EP�MQ�TZ	�B��  �у�_^[��]���������������������U���@SVW�EP�TZ	�Q��\  �Ѓ�_^[��]�������������������������U���\SVW�EP�MQ�U�R�TZ	�H��t  �҃����˝���M��[����E_^[��]��������������������������������U���PSVW�EP�M�Q�TZ	�B���  �у�P�M�i����M�话���E_^[��]�����������������U���PSVW�EP�M�Q�TZ	�B���  �у�P�M�����M��_����E_^[��]�����������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�E$P�M Q�UR�EP�MQ�UR�EP�MQ�TZ	�B���  �у� _^[��]�����������������������������U���@SVW�E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�TZ	�H���  �҃�$_^[��]��������������������������U���PSVWj �EP�MQ�UR�EP�M�Q�TZ	�B��t  �у�P�M�;����M�聛���E_^[��]�����������������������������������U���PSVW�EP�MQ�UR�EP�M�Q�TZ	�B���  �у�P�M�ȶ���M������E_^[��]���������������������U���@SVW�EP�TZ	�Q��8  �Ѓ�_^[��]�������������������������U���H  �B	3ŉE�SVW�E�E��E�P�MQh   ������R�t�����������Phȷ�TZ	�Q��4  �Ѓ��E�    _^[�M�3��������]���������������������������������U���DSVW�} 3��^�EP�MQ�UR�EP�	������E��}� |�E��9E�|/�}� }hз�lA	��P詚�����EE�@� �E���E��E�_^[��]�����������������������������������������U���PSVW�E�P�TZ	�Q��  �Ѓ�P�M�����M��S����E_^[��]���������������������U���PSVW�E�P�TZ	�Q��  �Ѓ�P�M轾���M������E_^[��]���������������������U���dSVW�n�����u�Vh���M�藢���EPh���M��L����EPh���M��;���j �E�PhicMC�M�Q�������M��v����M�����_^[��]��������������������������������U���dSVW�������u�M�����E�Xh!���M�������EPh!���M�豮��j �E�PhicMC�M�Q�f�����������P�M製���M��ܽ���M��I����E_^[��]�����������������������������������U���dSVW�>�����u�M�o����E�Xh����M��\����EPh����M�����j �E�PhicMC�M�Q�Ʒ�������O���P�M�����M��<����M�詘���E_^[��]�����������������������������������U���hSVW������u3��Rh#���M��Š���EPh#���M��z���j �E�PhicMC�M�Q�/��������W����E��M�諼���M������E�_^[��]����������������������������������U���hSVW������u3��Rhs���M��5����EPhs���M�����j �E�PhicMC�M�Q蟶������������E��M������M�舗���E�_^[��]����������������������������������U���@SVW�EP�MQ�UR�EP�MQ�UR�TZ	�H���  �҃�_^[��]����������������������U���@SVW�EP�MQ�UR�TZ	�H��@  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�EP�MQ�UR�TZ	�H���  �҃�_^[��]����������������������U���@SVW�E�8 t�E�Q�TZ	�B��D  �у��E�     _^[��]����������������������U���@SVW�EP�TZ	�Q��H  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q��L  �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�UR�TZ	�H��P  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H��T  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H��X  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H��\  �҃�_^[��]������������������U���@SVW�TZ	�H��d  ��_^[��]�����������������U���@SVW�E P�MQ�UR�EP�MQ�UR�EP�TZ	�Q��h  �Ѓ�_^[��]�����������������U���@SVW�EP�MQ�TZ	�B��l  �у�_^[��]���������������������U���@SVW�TZ	�H���  ��_^[��]�����������������U���TSVW�EP�M�Q�TZ	�B���  �у�P�M�����M�臓���E_^[��]�����������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�TZ	�B���  �у�_^[��]���������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H��l  �҃�_^[��]������������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���@SVW�EP�TZ	�Q���  �Ѓ�_^[��]�������������������������U���@SVW�EP�MQ�TZ	�B��$  �у�_^[��]���������������������U���@SVW�EP�TZ	�Q��(  �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q��,  �Ѓ�_^[��]�������������������������U���@SVW�TZ	�H��0  ��_^[��]�����������������U���@SVW�TZ	�H��<  ��_^[��]�����������������U���@SVW�EP�MQ�UR�EP�TZ	�Q���  �Ѓ�_^[��]�����������������������������U���@SVW�TZ	�H���  ��_^[��]�����������������U���@SVW�EP�MQ�UR�TZ	�H���  �҃�_^[��]������������������U���DSVWj �M�ܡ���E��}� t�E�P�N������E�P�ٟ����_^[��]����������������������U���@SVW�E$P�M Q�UR�EP�MQ�UR�EP�MQ�TZ	�B��  �у� _^[��]�����������������������������U���@SVW�TZ	�H��P  ��_^[��]�����������������U���@SVW�EP�MQ�UR�TZ	�H��`  �҃�_^[��]������������������U���DSVW�M��E���P蓫����_^[��]���������������U���@SVW�EP�TZ	���   ���   �Ѓ�_^[��]����������������������U���@SVW�EP�MQ�TZ	�Bd�HP�у�_^[��]������������������������U���@SVW�E�8 u��EP�TZ	�Qd�BT�Ѓ�_^[��]������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�Bh��у�_^[��]� �����������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�Bh���   �у�_^[��]� �������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Qh�B�Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�Hh�Q �҃�_^[��]� �������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�Bh���   �у�_^[��]� �������������������U���DSVW�M��EP�M�Q�TZ	�Bh���   �у�_^[��]� ���������������U���@SVW�TZ	�Hh�QX��_^[��]��������������������U���@SVW�E�8 u��EP�TZ	�Qh�B\�Ѓ�_^[��]������������������U���DSVW�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�TZ	�Bh�H`�у� _^[��]� ��������������������������U���DSVW�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�TZ	�Bh�Hd�у� _^[��]� ��������������������������U���DSVW�M��EP�MQ�U�R�TZ	�Hh�Qh�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�U�R�TZ	�Hh�Ql�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�U�R�TZ	�Hh�Qp�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Qh�Bt�Ѓ�_^[��]� ��������������������������U���@SVW�EP�MQ�UR�EP�MQ�TZ	�Bh���   �у�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�Bh�Hx�у�_^[��]� ������������������U���DSVW�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�TZ	�Bh���   �у� _^[��]� �����������������������U���DSVW�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�TZ	�Bh���   �у� _^[��]� �����������������������U���DSVW�M��E P�MQ�UR�EP�MQ�UR�EP�M�Q�TZ	�Bh���   �у� _^[��]� �����������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�Qh�B|�Ѓ�_^[��]� �������������������������U���DSVW�M��E P���E�$���E�$���E�$�M�Q�TZ	�Bh���   �у� _^[��]� ��������������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�Hh���   �҃�_^[��]� ����������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�Bh���   �у�_^[��]� �������������������U���@SVW�E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�TZ	�Hh���   �҃�$_^[��]��������������������������U���@SVW�E<P�M8Q�U4R�E0P�M,Q�U(R�E$P�M Q�UR�EP�MQ�UR�EP�MQ�TZ	�Bh���   �у�8_^[��]�������������������������������������U���@SVW�E@P�M<Q�U8R�E4P�M0Q�U,R�E(P�M$Q�U R�EP�MQ�UR�EP�MQ�UR�TZ	�Hh���   �҃�<_^[��]����������������������������������U���hSVW�M��M�������EP�M��?���P�M��z���j �M�Q�U�R�M�����M�襛���E�P�M�Þ���M������E_^[��]� �����������������������������U���DSVW�M��EP���E�$�M�Q�TZ	�Bh���   �у�_^[��]� ����������������������U���DSVW�M��EP���E�$�M�Q�TZ	�Bh���   �у�_^[��]� ����������������������U���DSVW�M��EP�MQ�U�R�TZ	�Hh���   �҃�_^[��]� ����������������������������U���DSVW�M��EP�MQ�U�R�TZ	�Hh���   �҃�_^[��]� ����������������������������U���\SVW�M��E(P�M$Q���E�$���E�$�UR�EP�M�Q�U�R�TZ	�Hh���   �҃�(�M���P�Q�P�Q�P�Q�P�Q�@�A�E_^[��]�$ ��������������������������������������U���\SVW�M��E$P���E�$���E�$�MQ�UR�E�P�M�Q�TZ	�Bh���   �у�$�U��
�H�J�H�J�H�J�H�J�@�B�E_^[��]�  �����������������������������������������U���DSVW�E�E��}�t��E�|Z	�E�xZ	�   _^[��]� ���������������������������U���PSVW�E�E��M����M��}��D  �U��$��F�   �3  ��Z	����Z	�=�Z	��   �EP������=�6  }
�������   �} u
�������   h(��pA	��PhH_	j�Z������E��}� t�M��(����E���E�    �M��tZ	�=tZ	 t�EP�tZ	�l����   �   �EP�MQ�:�������u����n�   �g�f����`��Z	����Z	uG���������=tZ	 t*�tZ	�E��M��M��}� tj�M������E���E�    �tZ	    �   ����_^[��]�vEBFIFlE�F"F��������������������������������������������������������������������������������������������������������U���@SVW�TZ	�HL���   ��_^[��]�����������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVW�TZ	�HL���_^[��]���������������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���DSVW�M��E�P�TZ	�QL���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�U�R�TZ	�HL���   �҃�_^[��]� ����������������������������U���HSVW�M��E�P�TZ	�QL���   �Ѓ��E��}� u j �EP�M�Q�TZ	�BL���   �у���M�豅��P�M�W���_^[��]� �������������������������U���DSVW�M��TZ	���   �M��BP��_^[��]�����������U���DSVW�M��E�P�TZ	�QL��(  �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�U�R�TZ	�HL��,  �҃�_^[��]� ����������������������������U���@SVW�TZ	�HL�Q��_^[��]��������������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���XSVW�M��EP�M�Q�U�R�TZ	�HL�Q�҃�P�M�ʓ���M��4|���E_^[��]� ���������������������������U���DSVW�M��EP�M�Q�TZ	�BL���   �у�_^[��]� ���������������U���DSVW�M��EP�MQ�U�R�TZ	�HL�Q�҃�_^[��]� ���������������U���DSVW�M��E�P�TZ	�QL�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QL�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QL�B�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QL�B �Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�M�Q�TZ	�BL��4  �у�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QL�B$�Ѓ�_^[��]� ��������������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�BL�H(�у�_^[��]� ����������������������U���DSVW�M��E�P�TZ	�QL�B,�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QL�B0�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�U�R�TZ	�HL��  �҃�_^[��]� ����������������������������U���DSVW�M��E�P�TZ	�QL���   �Ѓ�_^[��]����������������������U���XSVW�M��EP�M�Q�U�R�TZ	�HL��  �҃�P�M�����M��Qx���E_^[��]� ������������������������U���DSVW�M��E�P�TZ	�QL�B4�Ѓ�_^[��]�������������������������U���DSVW�M�j �E�P�TZ	�QL�B8�Ѓ�_^[��]�����������������������U���DSVW�M��EP�MQ�TZ	�BL�M����   ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�BL�M����   ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�BL�M����   ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�BL�M����   ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�BL�M����   ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�BL�M����   ��_^[��]� ���������������U���DSVW�M��EP�MQ�UR�EP�TZ	�QL�M���l  ��_^[��]� �����������������������U���DSVW�M��EP�TZ	�QL�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�QL�M����   ��_^[��]� �������������������U���DSVW�M��EP�TZ	�QL�M����   ��_^[��]� �������������������U���DSVW�M��EP�M�Q�TZ	�BL�H<�у�_^[��]� ������������������U���DSVW�M��E�P�TZ	�QL�B�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�U�R�TZ	�HL�Q@�҃�_^[��]� ���������������U���DSVW�M�j �EP�M�Q�TZ	�BL�HD�у�_^[��]� ����������������U���DSVW�M�j �EP�M�Q�TZ	�BL�HH�у�_^[��]� ����������������U���DSVW�M�j�EP�M�Q�TZ	�BL�HD�у�_^[��]� ����������������U���DSVW�M�j�EP�M�Q�TZ	�BL�HH�у�_^[��]� ����������������U���tSVW�M��M��o��h�  �M���|��P�M��	��j �E�P�M�Q�M��Qp��������E��M��*����U���t�E�    �M�胗���E���M������E��M��k����E�_^[��]������������������������������������������U���hSVW�M�j�M��8���h�  �M��|��P�M��W~��j�E�P�M�Q�M��x���M�肉���M�����_^[��]����������������������������U���hSVW�M��EP�M�膄��h�  �M��{��P�M���}��j�M�Q�U�R�M��x���M������M��x���_^[��]� �����������������������U���DSVW�M��E��     �E��@    �EP�M�Q�TZ	���   �H(�у��E�_^[��]� �������������������������U���hSVW�M��EP�M�趃��h�  �M���z��P�M��}��j�M�Q�U�R�M��@w���M��@����M�訕��_^[��]� �����������������������U���lSVW�M��M��.m��h�  �M��nz��P�M��|��j �E�P�M�Q�M���m��������E��M��ʇ���U���t�M������M��"����E��M���y��P�M�4����M������E_^[��]� ������������������������������������������������U���DSVW�M��E�P�TZ	���   �BL�Ѓ�_^[��]����������������������U���lSVW�M��M��.l��h�  �M��ny��P�M��{��j �E�P�M�Q�M���l��������E��M��ʆ���U���t�M������M��"����E��M���x��P�M�4����M������E_^[��]� ������������������������������������������������U���|SVW�M��M��nk��h�  �M��x��P�M���z��j �E�P�M�Q�M��1l��������E��M��
����U���t���]��M��e����E���M�貄���]��M��M����E�_^[��]��������������������������������������������U���DSVW�M��E�P�TZ	���   �B<�Ѓ�_^[��]����������������������U���tSVW�M��M��~j��h�  �M��w��P�M���y��j �E�P�M�Q�M��Ak��������E��M������U���t�E�    �M��s����E���M������E��M��[����E�_^[��]������������������������������������������U���lSVW�M��M���i��h�  �M��w��P�M��Iy��j �E�P�M�Q�M��j��������E��M��j����U���t�M豌���M�����E�,�M��>����M���P�Q�P�Q�@�A�M�蔑���E_^[��]� ������������������������������������������������U���DSVW�M��E�P�TZ	���   �BP�Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QL���   �Ѓ�_^[��]����������������������U���TSVW�M�j�EP�M�Q�U�R�TZ	�HL���   �҃��M���P�Q�P�Q�@�A�E_^[��]� ������������������������������U���TSVW�M�j �EP�M�Q�U�R�TZ	�HL���   �҃��M���P�Q�P�Q�@�A�E_^[��]� ������������������������������U���lSVW�M��M��g��h�  �M���t��P�M��w��j �E�P�M�Q�M��ah��������E��M��:����U���t�M聊���M�蒏���E�,�M������M���P�Q�P�Q�@�A�M��d����E_^[��]� ������������������������������������������������U���lSVW�M��M���f��h�  �M��t��P�M��Iv��j �E�P�M�Q�M��g��������E��M��j����U���t�M豉���M�����E�,�M��>����M���P�Q�P�Q�@�A�M�蔎���E_^[��]� ������������������������������������������������U���lSVW�M��M���e��h�  �M��>s��P�M��yu��j �E�P�M�Q�M���f��������E��M�蚀���U���t�M�����M������E�,�M��n����M���P�Q�P�Q�@�A�M��č���E_^[��]� ������������������������������������������������U���tSVW�M��M��.e��h�  �M��nr��P�M��t��j �E�P�M�Q�M���e��������E��M������U���t�E�    �M��#����E���M�跑���E��M������E�_^[��]������������������������������������������U���hSVW�M����E�$�M�����h�  �M��q��P�M���s��j�E�P�M�Q�M��n���M�����M�背��_^[��]� ����������������������������������U���DSVW�M��E��    �E��E�X�E�_^[��]� ����������������������U���hSVW�M��EP�M��H{��h�  �M���p��P�M��5s��j�M�Q�U�R�M��`m���M��`~���M��ȋ��_^[��]� �����������������������U���hSVW�M��EP�M��!x��h�  �M��p��P�M���r��j�M�Q�U�R�M���l���M���}���M��X���_^[��]� �����������������������U���DSVW�M��E��     �E��@    �EP�M�Q�TZ	���   �H,�у��E�_^[��]� �������������������������U���hSVW�M��EP�M��Qw��h�  �M��o��P�M���q��j�M�Q�U�R�M�� l���M�� }���M�舊��_^[��]� �����������������������U���hSVW�M��EP�M���v��h�  �M��Jo��P�M��q��j�M�Q�U�R�M��k���M��|���M�����_^[��]� �����������������������U���hSVW�M��EP�M��qv��h�  �M���n��P�M��q��j�M�Q�U�R�M��@k���M��@|���M�訉��_^[��]� �����������������������U���hSVW�M��EP�M��x��h�  �M��jn��P�M��p��j�M�Q�U�R�M���j���M���{���M��8���_^[��]� �����������������������U���lSVW�M��M��`��h�  �M���m��P�M��9p��j �E�P�M�Q�M��a��������E��M��Z{���U���t�M衃���M�貈���E�,�M��.����M���P�Q�P�Q�@�A�M�脈���E_^[��]� ������������������������������������������������U���tSVW�M��M���_��h�  �M��.m��P�M��io��j �E�P�M�Q�M��`��������E��M��z���U���t�E�    �M������E���M��w����E��M��ˇ���E�_^[��]������������������������������������������U���tSVW�M��M��>_��h�  �M��~l��P�M��n��j �E�P�M�Q�M��`��������E��M���y���U���t�E�    �M��3����E���M��ǋ���E��M������E�_^[��]������������������������������������������U���LSVW�M��M��K����E��}�t�}�t�}�t	�E�    ��E�   �E�_^[��]������������������������������U���DSVW�M��TZ	�PL�M����  ��_^[��]�����������U���hSVW�M��EP�M���r��h�  �M��:k��P�M��um��j�M�Q�U�R�M��g���M��x���M�����_^[��]� �����������������������U���hSVW�M��EP�M��u��h�  �M���j��P�M��m��j�M�Q�U�R�M��0g���M��0x���M�蘅��_^[��]� �����������������������U���hSVW�M��EP�M��t��h�  �M��Zj��P�M��l��h�   j�c����P�M�Q�U�R�M��f���M��w���M�����_^[��]� �������������������������U���@SVW�EE_^[��]�����������U���@SVW�EP�TZ	�Q���   �Ѓ�_^[��]�������������������������U���@SVW�EP�TZ	�Q���   �Ѓ�_^[��]�������������������������U���@SVW�TZ	�H���   ��_^[��]�����������������U���@SVW�TZ	�H���   ��_^[��]�����������������U���@SVW�E�Q�TZ	�B���   �у��E�     _^[��]��������������U���@SVW�EP�TZ	�Q���   �Ѓ�_^[��]�������������������������U���DSVW��r���E��}� u3��Oj �EP�MQ�UR�E�P�TZ	�Q��h  �Ѓ���u"�}� t�E�P�TZ	�Q@�B�Ѓ��E�    �E�_^[��]��������������������������������U���@SVWj �EPj �MQ�os����P�UR�EP�TZ	�Q��h  �Ѓ�_^[��]��������������������������������U���@SVW�EE_^[��]�����������U���@SVW�EP�MQ�UR�EP�TZ	�Q���   �Ѓ�_^[��]�����������������������������U���@SVW�E P�MQ�UR�EP�MQ�UR�EP�TZ	�Q���   �Ѓ�_^[��]�����������������U���DSVW�M��E�P�TZ	�QL�BL�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QL�BP�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QL���  �Ѓ�_^[��]� �����������������������U���DSVW�M��EP�M�Q�TZ	�BL��  �у�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�BL���   �у�_^[��]� ���������������U���DSVW�M��E�P�TZ	�QL�BX�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QL�B\�Ѓ�_^[��]� ��������������������������U���   SVW�M��bo���E��}� u3��k  �E�    �E�    �E�    �M��kW���M��;\���E��E��E؉EċEPh]  �M���i��j j �E�P�M��Z����u��   �M���U���E���E�E�}� ��   �M��p����E�E�E��E�Ph�   ��^������u�}�}� u�uj �M��T���E��}� u�`�E�P�M���a���E�P��w�����}� t�E�P�TZ	�Q@�B�Ѓ��E�    �l����E���t����M�� z���M��$Z����t����N�}� t�E�P�TZ	�Q@�B�Ѓ��E�    �E�P�ow����ǅx���    �M���y���M���Y����x���_^[��]� ��������������������������������������������������������������������������������������������������������U���DSVW�M��E��     �E��@    �E��@    �E��@    �E��@    �E��@    �E��@    �E�_^[��]��������������������������������������U���DSVW�M��EP�MQ�UR�TZ	���   �M��B��_^[��]� ����������������������������U���DSVW�M��EP�TZ	���   �M����   ��_^[��]� ����������������U���DSVW�M��EP�TZ	���   �M��B<��_^[��]� �������������������U���DSVW�M��E�P�TZ	�QL�B`�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QL�Bd�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�BL�Hh�у�_^[��]� ������������������U���DSVW�M��E�P�TZ	�QL��D  �Ѓ�_^[��]����������������������U���DSVW�M��E�P�TZ	�QL�Bl�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�BL���   �у�_^[��]� ���������������U���DSVW�M��E��M�H�E��M$�Hh`qh0qh qh�p�E��HQ�U R�EP�MQ���E�$�UR�E��HQ�U�R�TZ	�HL���   �҃�4_^[��]�  ���������������������������������������U���@SVW�E��M���_^[��]���������������������U���@SVW�EP�M��M�B��_^[��]����������������U���@SVW�EP�MQ�U��M�P��_^[��]������������U���@SVW�EP�MQ�UR�EP�M��M�B��_^[��]��������������������U���DSVW�M��E�P�TZ	�QL���   �Ѓ�_^[��]����������������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QL��   �Ѓ�_^[��]� �����������������������U���DSVW�M��EP�MQ�UR�EP�MQ�TZ	�BL�M���H  ��_^[��]� �������������������U���DSVW�M��TZ	�PL�M���L  ��_^[��]�����������U���DSVW�M��EP�TZ	�QL�M���P  ��_^[��]� �������������������U���DSVW�M��EP�TZ	�QL�M���T  ��_^[��]� �������������������U���DSVW�M��EP�MQ�TZ	�BL�M���p  ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�BL�M���t  ��_^[��]� ���������������U���DSVW�M��EP�MQ�UR�EP�MQ�U�R�TZ	�HL���   �҃�_^[��]� ����������������U���DSVW�M��EP�MQ�UR�E�P�TZ	�QL���   �Ѓ�_^[��]� �����������������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�BL��   �у�_^[��]� �������������������U���hSVW�M��3S���M��4r���} t�M��-R����u�E�   �M��?K���M���q���E��Kj�M��R��P�M�Z���M���Q���E��E�E�E�Ph=����U�����E��M���J���M��q���E�_^[��]����������������������������������������U���hSVW�M��sR���M��tq���} t�M��mQ����u�E�   �M��J���M��q���E��Kj�M��CQ��P�M��Y���M��2Q���E��E�E�E�Ph<���&U�����E��M��2J���M���p���E�_^[��]����������������������������������������U���@SVW�EP�MQ�UR�TZ	�HL���   �҃�_^[��]������������������U���@SVW�EP�MQ�TZ	�BL���   �у�_^[��]���������������������U���@SVW�EP�MQ�TZ	�BL���   �у�_^[��]���������������������U���@SVW�TZ	�HL��  ��_^[��]�����������������U���@SVW�TZ	�HL��@  ��_^[��]�����������������U���DSVW�M��EP�MQ�TZ	�BL�M����  ��_^[��]� ���������������U���DSVW�M��EP�MQ�TZ	�BL�M����  ��_^[��]� ���������������U���DSVW�M��EP�TZ	�QL�M����  ��_^[��]� �������������������U���DSVW�M��4S���M���E�_^[��]�����������������U���@SVW�TZ	���   ���   ��_^[��]��������������U���DSVW�M��E�P��k�����E��     _^[��]�������������������������U���DSVW�M��E�� _^[��]���������U���DSVW�M��и�]����z	�и�]����]����Au	����]�E�ش������$�y�����E���E��ش�X�M��e���E�_^[��]� ��������������������������������U���PSVW�M����]����Az	�E�   ��E�    ���]����Az	�E�   ��E�    �E�3�;E����M����E�$�1K����������$�Jx�����E�����E�$�K����������$� x�����E��X�E����X����Auh��tA	��P�L�����E����X�}� u�E�� ���M���M���c���E�_^[��]� ����������������������������������������������������������������������U���@SVW���E�$��n����_^[��]����������������U���DSVW�M��E��E�X�E����X����Auh��xA	��P�*K�����E����X_^[��]� ���������������������U���LSVW�M����]����Auh��|A	��P��J�������]�E�� �M���$�v�����M����A�$�]��v�����}����$�v�����U�����E�$�jv�����E��X�M��b��_^[��]� ��������������������������������������������������U���pSVW�M��E���� �$��H�����]�E����@�$�H�����]�����]�����At����]�����Au�E�����E����X�U  �H��]�����Auz�H��]�����Auj�E���V���E��E���V���E܃}� u�E�����E����X�8�E���}܉U؋E܉E��E؉E܃}� u��E��E��8�M���E��E��x�M��Y��   ���E��$���E��$�d�����=8��]����]�����Au.�E��M��]��E��M��]�E�� �MЋM���E��@�MЋM��Y���]�����Au���]�E����X���E��$���E��$�n�����]��E��]��E��]�����]�����A{ǋE�� �u�M���E��@�u�M��Y_^[��]������������������������������������������������������������������������������������������������������������������������U���@SVW�E�]����Au�E��E_^[��]������������U���@SVW���E�$���E�$�%n����_^[��]�����������������������U���@SVW�E��M�B��_^[��]��������������������U���@SVW�E��M�B��_^[��]��������������������U���DSVW�M��E�� X��E��@    h��E�Ph��h<��TZ	�QP��Ѓ��M��A�E�_^[��]�������������������������������U���DSVW�M�3�_^[��]������������U���@SVW�E��M�B��_^[��]��������������������U���DSVW�M��M��C���E��t�E�P�JL�����E�_^[��]� ����������������������������U���DSVW�M��E�� X��E��x u�E��HQ�TZ	�BP�H�у�_^[��]��������������������U���DSVW�M��E��x u3��"j �EP�MQ�U��BP�TZ	�QP�B�Ѓ�_^[��]� ����������������������������U���DSVW�M��E��x t�EP�M��QR�TZ	�HP�Q�҃�_^[��]� �����������������������U���DSVW�M��E��x t�EP�M��QR�TZ	�HP�Q�҃�_^[��]� �����������������������U���@SVW�TZ	�HP���   ��_^[��]�����������������U���@SVW�EP�TZ	�QP���   �Ѓ�_^[��]�������������������������U���@SVW�TZ	�HP�QP��_^[��]��������������������U���@SVW�EP�TZ	�QP�BT�Ѓ�_^[��]������������U���DSVW�M��E��     �E��@    �E�_^[��]������������������������U���DSVW�M��E��8 u�7�E��Q�TZ	�BP�HL�у��E��Q�TZ	�BP�H<�у��E��     _^[��]�����������������������������U���DSVW�M��EP�MQ�M��J��P�M��b��_^[��]� ������������������U���DSVW�M��E��@_^[��]��������U���HSVW�M��E��8 t*�E��Q�TZ	�BP�H<�у��E��     �E��@    �E��M�Hh��EPh��h<��MQ�UR�TZ	�HP�Q8�҃��M���E�    �	�E����E��E�;E}e�E��M���z u.�E��M���B   �E��M���BP�TZ	�QP�B�Ѓ��E�P�M��R�TZ	�HP�Q@�҃��M��U���A늋E�3Ƀ8 ����_^[��]� ��������������������������������������������������������������������U���LSVW�M��E�    �E�    �	�E���E�E��M�;H}a�E�P�M��R�TZ	�HP�Q@�҃��E��}� t!j �EPj�M�Q�TZ	�BP�H�у���u�E��Q�TZ	�BP�HL�у�3��닸   _^[��]� �������������������������������������������������U���DSVW�M��E��Q�TZ	�BP�HD�у�_^[��]�����������������������U���DSVW�M��E��Q�TZ	�BP�HH�у�_^[��]�����������������������U���DSVW�M��E��Q�TZ	�BP�HL�у�_^[��]�����������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���\SVW�M��E�P�M�Q�TZ	�BX��у��U��
�H�J�H�J�H�J�H�J�@�B�E_^[��]� ���������������������������U���\SVW�M��E�P�M�Q�TZ	�BX�H�у��U��
�H�J�H�J�H�J�H�J�@�B�E_^[��]� ��������������������������U���\SVW�M��E�P�M�Q�TZ	�BX�H�у��U��
�H�J�H�J�H�J�H�J�@�B�E_^[��]� ��������������������������U���   SVW�M��E�P��\���Q�TZ	�BX�H�у��   ���}�E_^[��]� �����������������������������U���DSVW�M��EP�M�Q�TZ	�BX�H�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�BX�H�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�BX�H�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�BX�H�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�BX�H$�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�BX�H �у�_^[��]� ������������������U���DSVW�M��EP�MQ�U�R�TZ	�HD�Q�҃�_^[��]� ���������������U���@SVWj �EP�TZ	�QD��Ѓ�_^[��]�����������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVW�EP�MQ�TZ	�BD��у�_^[��]�������������������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVWj �EP�TZ	�QD��Ѓ�_^[��]�����������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVW�EPh2  �TZ	�QD��Ѓ�_^[��]������������������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVW�EPhO  �TZ	�QD��Ѓ�_^[��]������������������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVW�EPh'  �TZ	�QD��Ѓ�_^[��]������������������������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVWj h�  �TZ	�HD��҃�_^[��]�����������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVWj h:  �TZ	�HD��҃�_^[��]�����������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���LSVW�M��M��H���E�    �E�    �E�Pj�M��J����u3���E�_^[��]�������������������������������U���DSVW�M��E��     �E��@    �E�_^[��]������������������������U���@SVWj h�F �TZ	�HD��҃�_^[��]�����������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���@SVWj h�_ �TZ	�HD��҃�_^[��]�����������U���@SVW�E�Q�TZ	�B@�H�у��E�     _^[��]�����������������U���LSVW�M��} u3��0�M���F���E�    �E�E��E�Pj�M��}H����u3���   _^[��]� ���������������������������������U���DSVW�M��E�P�TZ	�QD�B$�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B(�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�QD�B�Ѓ�_^[��]�������������������������U���DSVW�M��E��     �E��@    �E��@    �E��@    �E�_^[��]��������������������U���DSVW�M��M��2��_^[��]����������������������U���DSVW�M��E��     �E��@    �E��@    �E��@    �E�M�P;QuKjj�M��[����u�   �E���U���E���U�B�A�E���U�B�A�E��H�   �Tjj�M���Z����u�B�E���U���E���U�B�A�E���U�B�A�E���U�B�A�E��H�   �E�_^[��]� ��������������������������������������������������������������������U���DSVW�M��E��     �E��@    �E��@    �E��@    �EP�M��U���E�_^[��]� ���������������������U���DSVW�M��EP�M��^U���E�_^[��]� ������������U���DSVW�M��M��*0���} ��   hp���A	��P�M��Q�TZ	�B���   �у��U���E��8 u3��i�} tHhp���A	��
P�M��Q�TZ	�B���   �у��U��B�E��x u�E�P��?����3���E��M�H�E��M�H�   �3�_^[��]� ������������������������������������������������������U���DSVW�M��E�P�U?�����E���P�F?�����E��@    �E��@    _^[��]�������������������������������U���DSVW�M��M���.���} �	  �E�8 ��   �E�x ��   hp���A	��P�M�Q��R�TZ	�H���  �҃��M���E��8 u3��   �E�x tO�E�x tFhp���A	��
P�M�Q��R�TZ	�H���  �҃��M��A�E��x u�M��.��3��^�E��M�Q�P�E��M�Q�P�E��HQ�U��P�M�R�BS�����E��x t�E��HQ�U��BP�M�QR�S�����   _^[��]� �������������������������������������������������������������������������������������������U���DSVW�M��M��:-���} �D  �} �:  hp���A	��P�M��Q�TZ	�B���  �у��U���E��8 u3��  �} tX�} tRhp���A	��
P�M��Q�TZ	�B���  �у��U��B�E��x u�M��,��3��   �E��M�H�P�E��@   hp���A	��P�M��Q��R�TZ	�H���  �҃��M��A�E��x u�M��?,��3��T�E��M�H�E��HQ�U��P�MQ�~Q�����} t�E��HQ�U��BP�MQ�^Q������E��H�U��   _^[��]� ������������������������������������������������������������������������������������������������U���DSVW�M��E��     �E��@    �E��@    �E��@    _^[��]�����������������������U����  SVW�M����]��E�    j �M���4��j �M���4��j �M���4���E��H�U�<�}���E  �} ��  �M��VG��j ��t����4���E���k�U��EԋJ�M؋B�E܋J�M��B�E�J�M�E�P�M���Bk�EP��<���Q��@�������t����H��x����P��|����H�M��P�U��@�E��E�   �	�E����E��E��H�U�;��   �E�P�M���E���k�MQ��T���R�@������M��P�U��H�MċP�UȋH�M̋P�UЍE�P��t���Q��l���R��7����P�M��0���E���t����M���x����Uĉ�|����EȉE��M̉M��UЉU��I��������$��������6���E��������������P�������H�������P�������H�������P�E�P������Q�?�����U��H��
�H�J�H�J�H�J�H�J�@�B���E��$�&���E��$ݝ4����&����ܝ4���������   ���E��$�^&���E��$ݝ4����M&����ܝ4���������   �E��HP�����$�����$�����$�������~4��P������Q�t6�����U����
�H�J�H�J�H�J�H�J�@�B�E��P�M��HQ������R�/6�����M��0���P�Q�P�Q�P�Q�P�Q�@�A�  ���E��$�%���E��$ݝ4����n%����ܝ4���������   �����$�����$�����$�������3��P�E��HP�����Q�5�����U����
�H�J�H�J�H�J�H�J�@�B�E��P�M��HQ��,���R�P5�����M��0���P�Q�P�Q�P�Q�P�Q�@�A�   �����$�����$�����$��D�����2��P�E��HP��\���Q��4�����U��0��
�H�J�H�J�H�J�H�J�@�B�E��HP�M��0Q��t���R�4�����M�����P�Q�P�Q�P�Q�P�Q�@�A�EP������Q�p7�����   ���}��E�    �	�E����E��E�;E}�E��H�U��E���E��ۋE���U��k�EP�MQ������R�<������MԋP�U؋H�M܋P�U��H�M�P�U�E���U�D�k�EP�MQ�����R�O<������M��P�U��H�MċP�UȋH�M̋P�U��E�    �	�E����E��E��H�U�E�;���   �E����M��I�u��<�U�E����k�UR�EP�����Q��;������U��H�M��P�U��H�M��P�U��@�E��E�P�M�Q�U�R�U  ���E��]�E��EԋM��M؋UĉU܋EȉE��M̉M�UЉU�E��E��M��M��U��UċE��EȋM��M̋U��U�� ����E�_^[��]� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���DSVW�M��E��M� ��U���E��M�@�A�U��Z�E��M�@�A�U��Z�E�_^[��]� ���������������������U���@SVW�E�M�@(�	�U�B�E�M�@@�I���U�E�BX�H�����$�M�U�A �
�E�@�M�U�A8�J���E�M�@P�I�����$�U�E�B��M��U�E�B0�H���M�U�AH�J�����$�M��-���E_^[��]����������������������������������������������U���@SVW�E�M�@�a�U�
�E�M�@�a�U�
���E�M�@�a�U�
��_^[��]��������������������������U���DSVWj�0   ���E��}� u3���E��H��_^[��]������������������U���@SVWh�Z	�EPh_� �>L����_^[��]�����������U���HSVW�E�8 u�5j�������E��}� u� �E��M��E�P�M��Q�҃��E�     _^[��]����������������������������������U���HSVW�M�j�M������E��}� t	�E��x u3���EP�U��M��B��_^[��]� ����������������������������U���HSVW�M�j��������E��}� t	�E��x u3���EP�U��M��B��_^[��]� ����������������������������U���HSVW�M�j�������E��}� t	�E��x u3���EP�MQ�UR�E��M��P��_^[��]� ��������������������U���HSVW�M�j�-������E��}� t	�E��x u3���EP�U��M��B��_^[��]� ����������������������������U���HSVW�M�j ��������E��}� t	�E��x  u3���EP�U��M��B ��_^[��]� ����������������������������U���HSVW�M�j$�m������E��}� t	�E��x$ u2���EP�U��M��B$��_^[��]� ����������������������������U���HSVW�M�j(�������E��}� t	�E��x( u3���E��M��P(��_^[��]�������������������U���HSVW�M�j,�������E��}� t	�E��x, u3���E��M��P,��_^[��]�������������������U���HSVW�M�j0�m������E��}� t	�E��x0 u3���EP�U��M��B0��_^[��]� ����������������������������U���HSVW�M�j4�������E��}� t	�E��x4 u�����EP�MQ�U��M��B4��_^[��]� �����������������������U���HSVW�M�j8�������E��}� t	�E��x8 u3���E��M��P8��_^[��]�������������������U���HSVW�M�j<�]������E��}� t	�E��x< u��EP�U��M��B<��_^[��]� ������������������������������U���HSVW�M�j@��������E��}� t	�E��x@ u��EP�U��M��B@��_^[��]� ������������������������������U���HSVW�M�jD�������E��}� t	�E��xD u3���EP�U��M��BD��_^[��]� ����������������������������U���HSVW�M�jH�=������E��}� t	�E��xH u��EP�U��M��BH��_^[��]� ������������������������������U���HSVW�M�jL��������E��}� t	�E��xL u3���E��M��PL��_^[��]�������������������U���HSVW�M�jP�������E��}� t	�E��xP u3���E��M��PP��_^[��]�������������������U���HSVW�M�jT�=������E��}� t	�E��xT u��E��M��PT��_^[��]���������������������U���HSVW�M�jX��������E��}� t	�E��xX u��E��M��PX��_^[��]���������������������U���HSVW�M�j\�������E��}� t	�E��x\ u��E��M��P\��_^[��]���������������������U���HSVW�M�j`�M������E��}� t	�E��x` u3���EP�MQ�U��M��B`��_^[��]� ������������������������U���HSVW�M�jd��������E��}� t	�E��xd u3���EP�MQ�U��M��Bd��_^[��]� ������������������������U���HSVW�M�jh�������E��}� t	�E��xh u��EP�MQ�UR�EP�MQ�U��M��Bh��_^[��]� ������������������������������U���HSVW�M�jl�������E��}� t	�E��xl u3���EP�MQ�UR�E��M��Pl��_^[��]� ��������������������U���HSVW�M�jp�������E��}� t	�E��xp u3���EP�MQ�U��M��Bp��_^[��]� ������������������������U���HSVW�M�jt�]������E��}� t	�E��xt u3���EP�MQ�U��M��Bt��_^[��]� ������������������������U���HSVW�M�jx��������E��}� t	�E��xx u3���EP�MQ�U��M��Bx��_^[��]� ������������������������U���HSVW�M�j|�������E��}� t	�E��x| u3���EP�U��M��B|��_^[��]� ����������������������������U���HSVW�M�h�   �:������E��}� t�E����    u3���EP�MQ�U��M����   ��_^[��]� �������������������������������U���HSVW�M�h�   ��������E��}� t�E����    u����&�EP�MQ�UR�EP�MQ�UR�E��M����   ��_^[��]� ������������������������������U���HSVW�M�h�   �J������E��}� t�E����    u����&�EP�MQ�UR�EP�MQ�UR�E��M����   ��_^[��]� ������������������������������U���HSVW�M�h�   ��������E��}� t�E����    u3���EP�MQ�UR�EP�U��M����   ��_^[��]� �����������������������U���HSVW�M�h�   �Z������E��}� t�E����    u3���EP�U��M����   ��_^[��]� �������������������U���HSVW�M�h�   ��������E��}� t�E����    u��EP�U��M����   ��_^[��]� ���������������������U���HSVW�M�h�   �������E��}� t�E����    u3���EP�MQ�U��M����   ��_^[��]� �������������������������������U���HSVW�M�h�   �*������E��}� t�E����    u3���EP�MQ�UR�E��M����   ��_^[��]� ���������������������������U����   SVW�M��M��@/���E�    �	�E����E��E��M�;H�  �E���U����97����u�ҋE���U�����%����E�E܋E܋M܋P;Qul�E܋k�MQ�U܋Bk�EP�����Q�(����P�U܋k�EP�M܋Qk�UR��$���P�(����P��<���Q� ����P�M������h�E܋k�MQ�U܋Bk�EP��T���Q�M(����P�U܋Bk�EP�M܋Qk�UR��l���P�#(����P�M�Q�����P�M����������E�P�MQ��'�����E_^[��]� ������������������������������������������������������������������������������������������������������U���   SVW�M��M��3���E�    �	�E����E��E��M�;H��   �E���U����i5����u�ҋE���U����$����E�E��E��k�MQ�M��7���E��Hk�MQ�M��7���E��Hk�MQ�M��7���E��M��P;Qt�E��Hk�MQ�M��n7���S����EP�MQ�M��k��_^[��]� ����������������������������������������������������������U���tSVW�M��M��S,���M����H,��������$�M�� ���E��M���U��P�M��H�U��P�M��H�U��P������$�M������E����M���U��P�M��H�U��P�M��H�U��P�E��@0    �E�_^[��]�������������������������������������������������������U���DSVW�M��E��x0 ��   �E�M�������Au
�E��M���E�M��A�X����Au�E��M�A�X�E�M��A�X����Au�E��M�A�X�E�M��A�����z�E��M��X�E�M��A �X����z�E��M�A�X �E�M��A(�X����z�E��M�A�X(�`�E�M������P�Q�P�Q�P�Q�P�Q�@�A�M����U����A�B�A�B�A�B�A�B�I�J�E��@0   _^[��]� ����������������������������������������������������������������������������������������U���   SVW�M��E��x0 ��   ������$�E���P�M�Q��\���R������P��t���P��	�����M���P�Q�P�Q�P�Q�P�Q�@�A�EP�M���Q�U�R�h#�����M���P�Q�P�Q�P�Q�P�Q�@�A�^�����$�M�����E�M���U��P�M��H�U��P�M��H�U��P�E�M���P�Q�P�Q�P�Q�P�Q�@�A_^[��]� ������������������������������������������������������������������������������������U���@SVW�E�@�M���$�M�A�M���$�U��M���$�M�����E_^[��]��������������������������U���LSVW�M��E�    �E��x|�E��8 u3��?�E�    �	�E���E�E��M�;H}�E���U���~����t	�E����E��͋E�_^[��]�����������������������������������U���DSVW�M��E�� %    _^[��]��������������������U���HSVW�M��E�E��	�E����E��E��M�;H}!�E���U���������t�E�+E����˃��_^[��]� ���������������������������U���HSVW�M��} |�E��8 u����<�E�    �	�E����E��E��M�;H}�E���U������;Eu�E���Ѓ��_^[��]� ����������������������������U���LSVW�M��E� �E�    �	�E���E�E��M�;H}3�E���U��� ��;Eu�]��E���U��������؈]���E���_^[��]� ���������������������������������U���HSVW�M��M�����E��}��u3��
�   �M���_^[��]���������������U���DSVW�M��E����   @t�����E�� %���3ҹ   ���_^[��]�����������������������U���LSVW�M��E�    �E�    �	�E���E�E��M�;H} �E���U���W�����t	�E����E��̋E�_^[��]�����������������������U���LSVW�M��E�    �E�    �	�E���E�E��M�;H}�E���U����,����t	�E����E��͋E�_^[��]������������������������U���PSVW�M��E�    �	�E����E��E��M�;H}�E���U���%����M���M������E�    �	�E����E��E��M�;H}{�E���U���%   �ud�E���U��������E��E����E��	�E���E�E��M�;H}2�E���U�����;E�u�E���U��   ��M���M����q���_^[��]������������������������������������������������������������U���LSVW�M��M��)����E�E��M��r���E��E����E��}�wz�M��$�<��E� ����E� ����\�E�M����E�M��Q��E�E�M��Q��E�M��Q��-�E�M��Q��E�M��Q���E�M��Q��E�M���_^[��]� ��������������������������������������������������������������������������U���LSVW�M��M�����E��M��h���E�E;E�t	�}���u�E;E�t	�}���u�^�}���t�E�E�}���t�E�E��}��t�E��M���E����   �ыE����E���   @�M����   �M��_^[��]� ���������������������������������������������������U���@SVW�E��P�MQ�UR������_^[��]����������U���@SVW�TZ	�H\���_^[��]���������������������U���@SVW�E�Q�TZ	�B\�H�у��E�     _^[��]�����������������U���DSVW�M��E�P�TZ	�Q\�B�Ѓ�_^[��]�������������������������U���DSVW�M��E�P�TZ	�Q\�B�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�B\�H�у�_^[��]� ������������������U���DSVW�M��EP�MQ�U�R�TZ	�H\�Q�҃�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�B\�H�у�_^[��]� ������������������U���DSVW�M��E�P�TZ	�Q\�B�Ѓ�_^[��]�������������������������U���DSVW�M��EP�M�Q�TZ	�B\�H �у�_^[��]� ������������������U���DSVW�M��EP�MQ�U�R�TZ	�H\�Q$�҃�_^[��]� ���������������U���DSVW�M��EP�MQ�UR�EP�M�Q�TZ	�B\�H`�у�_^[��]� ����������������������U���DSVW�M��EP�M�Q�TZ	�B\�H0�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�B\�H@�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�B\�HD�у�_^[��]� ������������������U���DSVW�M��EP�M�Q�TZ	�B\�HH�у�_^[��]� ������������������U���DSVW�M��E�P�TZ	�Q\�B4�Ѓ�_^[��]�������������������������U���DSVW�M��EP�MQ�U�R�TZ	�H\�Q8�҃�_^[��]� ���������������U���DSVW�M��EP�M�Q�TZ	�B\�H<�у�_^[��]� ������������������U���TSVW�M�j �M�����M��z���E�E�P�M����E�    �	�E����E��E�;E�}3�E�P�M�Qh����U�R�M���+���E�P�M�q���E�P�M�e���_^[��]� ���������������������������������������������U���XSVW�M��E�P�M�(����}� |o�M������E�P�M�����}� tU�E�    �	�E���E�E�;E�};�E�P�M������E�P�M������	�E���E�E�;E��E�P�M������봸   _^[��]� �����������������������������������������������������U���H  �B	3ŉE�SVWh    ��Z	P��������t
������Z	jjj�#����P�#����P�EP��Z	Q������P�}�������u��   �E������������P�MQh�  ������R�>����j�EP�>�������th��������j�EP��������th�������������P�����h   @�EP���������t�EP�MQ�3  ��h    �EP���������uh ��j����ǅ����    _^[�M�3���'����]������������������������������������������������������������������������������������U���@SVW�E#E_^[��]�����������U���@SVWh    jjj��!����P��!����P��!����_^[��]����������������������������U���@SVW�EPhȷ�����_^[��]����������������U���  �B	3ŉE�SVW�E�P��   ���E�P�   ���E��E�Ph0�j?�M�Q������EP�MQ�U�Rh �h�  ������P�! ����������P������_^[�M�3��e&����]������������������������������������U���@SVW�EP�C�����_^[��]���������������������U���@SVW�EP�����_^[��]���������������������U���HSVW�} 3��   �E�E��E�P�MQ�UR�EP�@�����E��}� |�E�;E|l�}� }Sh@���A	��	PhH�h@�hH������P�	����Ph   @j������P�b������Z	��t̋EE�@� �E���E��E�    �E�_^[��]���������������������������������������������������������������U���@SVW�̑	�����_^[��]���������������������U���@SVW�E�M��E�M�H�EPj�MQ�j����_^[��]��������������U���@SVW�   _^[��]������������U���HSVW�} t�E�8 t�E� �Pj�EP��������E��}� u3��5�M������E��}� u3�� �} t�E�M���E��M;H~3���E�_^[��]��������������������������������������������U���LSVW�M��EP�TZ	�Q�M��Bd�ЉE��}� u3��ah����A	��P�M���Q�TZ	�B���   �у��E�}� u3��+�EP�M���Q�U�R�TZ	�P�M��Bh�ЋE�E��  �E�_^[��]� ����������������������������������������U���@SVWj h�  h�Z	�M�����Z	_^[��]������������������������U���@SVWj h�  h�Z	�M������Z	_^[��]������������������������U���@SVWh� �M�o����tj h�  h�Z	�M�p��������h�h�Z	��������Z	_^[��]����������������������������U���DSVW�M��EP�TZ	���   �M��B��_^[��]� �������������������U���PSVWj h�  h�Z	�E�P�M������������M�������Z	_^[��]���������������������U���PSVWj h�  h�Z	�E�P�M����������M��������Z	_^[��]���������������������U���`�B	3ŉE�SVW�E�E��E�    �E��D�0�M���M�E��D�x�M���M��E�   �	�E���E�}� |I�E��M������E��E��
}�E��0�M�D�U���U���E��7�M�D�U���U�먋E��D� j �E�P�M����E_^[�M�3��U ����]����������������������������������������������������U����   SVW�} ��   �}   @��   j h,���@������Pj0j jj �E�U��������8�����<���߭8����5 ����$��P���P�9�����P�MQ�J������P���������@��������E�F  �  �} ��   �}   ��   j h���`���� ��Pj0j jj �E�U�
�D�����8�����<���߭8����5 ����$��p���P������P�MQ�������p����u�����`����j����E�   �f�} |`	�}   vUj h��M��p��Pj0j jj �m�5 ����$�E�P�*�����P�MQ�;�����M������M�������E�@j h��M����P�EP�M�Q�K����P�UR�������M�������M������E_^[��]�������������������������������������������������������������������������������������������������������������������������������U���PSVW�E P�MQ�UR�EP���E�$�M�Q�TZ	�B�H$�у�P�M����M�������E_^[��]��������������������̋�U���uQ���YY]� ����̋�Q�4��r���Y����̋�U��V��������EtV�r���Y��^]� �������̋�U���uQ�����YY]� ����̋�Q�X��Y��̋�U��E��	Q��	P�������Y�Y@]� �������̋�U��E��	Q��	P������Y�Y��]� �������̋�U��E��	Q��	P�p���YY3Ʌ�����]� ��������̍AË�� 4�� �̋�� ��� B	�$B	��(B	��,B	���0B	���4B	�8B	o��<B	���@B	}��DB	 �������������������������̋�U��M�L_	�L_	]�����̋�U������} t������]���������������̃=��	 t-U�������$�,$�Ã=��	 t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$��������������������������������������������jh�'	�
���E��uz�=�����u3��8  ������u�������
���ؑ	�̄	�q���T_	�����y� ����������x �Z����xj ����Y��u�P_	��   ������3�;�u[9=P_	~��P_	�}�9=�_	u�����9}u�V���� ���
����E������   �   3�9}u�=PB	�t� ����j��uY�T���h  j����YY��;�����V�5PB	�5|_	�ԑ	�Ѕ�tWV���YY�Б	��N��V�?��Y�������uW�L���Y3�@����� �����������������������������������������������������������������������������������������jh�'	��������]3�@�E��u9P_	��   �e� ;�t��u.�@���tWVS�ЉE�}� ��   WVS�����E����   WVS������E��u$��u WPS����Wj S����@���tWj S�Ѕ�t��u&WVS�����u!E�}� t�@���tWVS�ЉE��E������E���E��	PQ�6���YYËe��E�����3�����������������������������������������������������������������̋�U��}u�����u�M�U����Y]� �������̋�U��QSV�5ԑ	W�5��	���5��	�؉]��֋�;���   ��+��G��ruS�4����؍GY;�sH�   ;�s���;�rP�u��O��YY��u�C;�r>P�u��9��YY��t/��P�4��ܑ	���	�u�=ܑ	�׉��V�ף��	�E�3�_^[����������������������������������������������̋�Vjj ����YY��V�ܑ	���	���	��ujX^Ã& 3�^�������������jh(	�J������e� �u�����Y�E��E������	   �E�������)�����������������̋�U���u���������YH]��������������̋T$�L$��ti3��D$��u���   r�=��	 t�����W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$��������������������������������������̃=<�	 ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�y[  ��=<�	 t2���\$�D$%�  =�  u�<$f�$f��f���d$u�h������$�����   ��ÍT$�>���R��<$tPf�<$t�-8�������z�=L_	 ����   ��A	�S���-:���������z��������.������� u�|$ u����-���   �=L_	 �����   ��A	�[��Z���������������������������������������������������������������������������������������̃=<�	 ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�`  ��=<�	 t2���\$�D$%�  =�  u�<$f�$f��f���d$u�D������$�[���   ��ÍT$����R��<$tmf�<$t�g��=  �?s+��������������=L_	 �����   ��A	����w:�D$��%�� D$u)��   ����-��t������������ u�|$ u����-���   �=L_	 �)���   ��A	���Z������������������������������������������������������������������������������������������̃��$�6
���   ��ÍT$����R��<$�D$tQf�<$t�>
���   �u���=L_	 �r���   � B	����  �u,��� u%�|$ u�������"��� u�|$ u�%   �t����-���   �=L_	 ����   � B	���Z����������������������������������������������̋�U��=a	 u����j����h�   �j���YY�E��u@Pj �5a	���	]���������������̋�U��S�]���woVW�=a	 u���j�>���h�   ����YY��t���3�@Pj �5a	���	����u&j^9xh	tS����Y��u������0����0��_^�S�����Y����    3�[]�������������������������������������̋�U��} t-�uj �5a	��	��uV�A������	P�J���Y�^]������������������������U��WV�u�M�}�����;�v;���  ���   r�=��	 tWV����;�^_u�7�����   u������r)��$�@��Ǻ   ��r����$�T��$�P���$����d�����#ъ��F�G�F���G������r���$�@��I #ъ��F���G������r���$�@��#ъ���������r���$�@��I 7�$����������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�@���P�X�d�x��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$����I �Ǻ   ��r��+��$����$�������<��F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I �����������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̃=<�	 ������\$�D$%�  =�  u�<$f�$f��f���d$����� �~D$f(`�f(�f(�fs�4f~�fT��f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�7������D$��~D$f��f(�f��=�  |!=2  �fTP��\�f�L$�D$����f���fV��fTp�f�\$�D$��������������������������������������������������������������������������������U��WV�u�M�}�����;�v;���  ���   r�=��	 tWV����;�^_u������   u������r)��$����Ǻ   ��r����$���$� ���$�����@�d�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I �����������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$����� ���(��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�<��I �Ǻ   ��r��+��$����$�����������F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I @�H�P�X�`�h�p����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+������������������������������������;B	u��������̋�U��QQ��VW�]����  Vh?  ����YY�M����  #�f;�uh�EQQ�$����HYYtJHt9H�EWt!������\$�E�$jj�������HQQ�$j�{������7VW�����E���'VW�����E��E%����E��EVW�E��o����E�YY_^�������������������������������������������������������̺�����������������������z�������������5Dl	�ԑ	��t��j�v���jj ��������������������̋�U��V�5Dl	�ԑ	�u���ܑ	�Dl	��^]�����������5Dl	�ԑ	���̋�U��� �e� Wj3�Y�}��9Eu�����    �[ ������x�MV�u��t��u�����    �7 ������S�����E�;�w�M��u�E��u�E�B   �u�u�P�u��Q���������t�M�x�E��  ��E�Pj ����YY��^_��������������������������������������������̋�U���uj �u�u�u������]�������̋�U��} t�u�u�u�u�u����]��������̋�U��EV���F ��uc�����F�Hl��Hh�N�;�N	t�L	�Hpu�������F;J	t�F�L	�Hpu�����F�F�@pu�Hp�F�
���@�F��^]� ��������������������������������̀y t�A�`p����̋�Ë�U��E��t�M���]�����̋�U��E��t���8��  uP����Y]��������̋�U���SVW�u�M�3������E苸�   �]��u��t������4��E�������E��}�YY�M��\rՍCP������Y�u���td�e� �E��:�4��E�F+ƍDPV��������uTV������E��:�t��E�F+ƍDPV�}�������u*V������E��}�Yr�� �}� _^[t�E��`p��E���3�PPPPP���������������������������������������������������������������j ����Y��̋�U���SVW�u�M�3��z����E䋸�   �w8�u��E�   �v0������6�E�������u�YY�M�Ã��M��\�u�uՍCP�������Y�u���tb�e� ��h�E��:�w�F+ƍDPV�p�������uRV������E��:�7F+ƍDPV�K�������u-V�Z�����E����}�Yr�� �}� _^[t�E�`p��E���3�PPPPP�a����������������������������������������������������������������j �����Y��̋�U���$SVW�u�M�3��C����E܋��   �}��]��t������4��E�������E��}�YY�M�|rՍF8�E��E�   �]��s0�x����3�E��n����E�YY�M���M�|u����   �O������   ���B������   Ǎ|�1������   �|�"������   �|������e  P�E��(����؃�����  hd  VS��d  ������e� �F�]���)u��E�E��<��E��p��+�E�PW��������uTW�����M��|�E�<�0��+�E�PW�q�������u*W�����E��E��}�Y�|r��e� �Ch�E�F8�E��3�PPPPP�����E�M��<�0��+�E�PW��������u�W�*����|�E�8�E��p0��+�E�PW���������u�W� ����E��E��E��}�Y�|r���+�E����   ���   PW���������i���W�����|��+�E����   ���   PW���������:���W�����|��+�E����   ���   PW�V�����������W�a����|��+�E����   ���   PW�'������������W�2����D��+�M����   ���   QP���������������}� t�E�`p�_^��[��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������j �)���Y��̃8 V��tW���t�9��F��8 u�_^��������̃>�Svj
�[����0�A����~��w��I���I�@;�r�[�������������̋�U��QSV��3҉U�9Ut5�9�7vj
�[����0�F�	���~��w��7N���N�@;�r��.;1s(N�V��tj
�[�����0�E��N���u�E�)��^[�������������������������������̋�U��QS��V�uW�ً���Y��  �{  ��I��   ��   ���v  ��	�m  ��tj��tEHt"���t  �F���Y  ���P  ��  �v���@  ���7  �U�T�h�  �v���   ���  �U�T���  �� %����  �v����  ����  �ƙjY����uQX���Q  ��M��   jY+�twHHt,HHtH��  �i  �F����  ;���  ��t�H���F����  ;��  �ȋF���r  =m  �g  ;�}3��j�^��;��x���@�r�������A  ��;�8  �Z����F���(  ��;������F=�����  =�  �  �jdY���u��j��k�d��t��m�  �  ��Z�%  ����   H��   HtUHt*����   �v����   ��m  ��   �u�Fj��v����   ����   ���ujZ� ���Y�c  �} �uSWVt<j�u�C  ����tc�; t^��  ���uSWVj�u�  �����  �8j �v��x���U�T�8��   �v��x��~������    ����3���   �U����   �v��x׃�ҍF�I�����p��   ��t]Ht@Ht$Hu������8�����3�9F ���E��Ë]����~�F��x��u�jdY���ˋ�������} �uSWVtj�)���j �"����F���T������K����u3�B������v���5������,����U�����   ����   �Ë��L���3�@_^[�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���0�B	3ŉE��E�M�� �E��ES�]V�u�E؋EW�E�tIt���   ����   ����   ���   ��  �}��	u��	�EԋEعl  fHf�M�f�HfAf�M�f�Hf�M�f�Hf�M�f�Hf� f�E�3�PPWf�M��M�QPf�E��E����   �UԉEЅ��  ��=   �X����ą�t� ��  �P����Y��t	� ��  ���E����   �uЉE�PW�E�P�E�j ���   �U�H��~�}�; v����G�H����u�����Y3�@�e�_^[�M�3�������3�9t�U��AB8t��M��ȃ�d�|  �H  ��'��   ��A��   ��Ht{��MtL��a��   �u�Q�(���YY��t�;v� ��  ����G�����G�����w����]�����HtHtHt
Hu��B�/  �b�(  �E�   �m�  ��HtHt	��E�   �H�  h(�W�7���YY��u���h$�W�!���YY��u���}�p��  ����p������������; �]���<'tB�u���P�J���YY��t�;v� ��  ����G�����G����u�����G������HtHtHtH������A�K  �a�D  �E�   �d�6  ����h�  ����   ����   Ht%��������B�HtHH�x����Y��   �y��   �E؃x�E����   ����   ����   �; v{��u�P�g���YY��t�;v� ��   ����G�������   �; ��   �u���P�#���YY��t�;v� ��   ����G�����G����u��b��HtHt�����E�   �S�.��HtHt�����E�   �M���HtHt�����E�   �I�u���u܋��u��u���������t�}�����3�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� �ES�u3ۍM��]��E��s����E;�u#�]����    ����8]�t�E�`p�3��@  W�};�u#�2����    �����8]�t�E�`p�3��  V�u�;���   �E;�u	�E����   �E�}�;���   �:�ty<%tA�M���QP����YY��t3�A9M�v�F8tp��U�
�E�M�����M��EF�M��/9]tyF3��>#u@FP�u�E��u�M�P��U���������tBF9]�w�9]�v�E�+}���8]�tT�M�ap��K�M��E��9]�u 9]�w�5���� "   �9]�v��E�   �������    ����8]�t�E�`p�3�^_[����������������������������������������������������������������������������������������������������̋�U���uj �u�u�u�u�:�����]��������̋�U��j j �u�u�u�u������]�������̋�U��j �u�u�u�u�u������]��������̋�U���V�uW3��}��}�}�;�u����j^�0�������TSj$h�   V�i����]��;�u�����j^�0�|����(�C�;�|;�r��|���o@�v����j^�0��[_^�������E�P����Y����  �E�P�����Y����  �E�P�r���Y����  �K�;��|j���� v`�E��+��E�P�V�}�M�����YY��u�9E��;  V����Y���,  �E��)E�E�PU�V�����YY���Y����F    �  SV�����YY���<���9E�t,V�p���Y��t!�E�E��F    ��ȋ�U�����+�]������E��ڙ+��j j<SW�������y��<��ĉ���j j<SW�h������F�ڙj �j<�SW������F��y��<��ĉF���j j<SW�3������F�ڙj �j�SW�����F��y�����F���j jSW������ȅ�|+��t�F�j�_��N�VN3��D������|��s�F�D�j_��N�F�V��ҁ�m  N���N�F�F   �WWWWW�d���������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��V���������t�uV�}������Y��Y#�^]���������̋�U��QQ�E�P���	�E��M�j  ��*h��� ��!Nb�QP������|=�o@�v����ЋM��t��Q������������������������������������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_������������������������������������������������������������������������̀�@s�� s����Ë���������������������jh8(	����j�f���Y�e� �u�N��t/�l_	�h_	�E��t9u,�H�JP�o���Y�v�f���Y�f �E������
   �"���Ë���j�����Y�����������������������������jhX(	�%����}3�9_��   h (  h��h~�S�G	PS�B������E�;�u3��   P����Y���N�E�<0 u�0;�w�Nj����Y�]�9_uVj����Y�؅�tH��V�p���Y�G��t0�u�VP�8�����3�;�u�G��E�H�K�X�QQQQQ�h���S�_���Y�u��V���Y�E������   �G����Ë}j�����Y�������������������������������������������������������������jhx(	�����j����Y�e� �u�N��t/�l_	�h_	�E��t9u,�H�JP����Y�v����Y�f �E������
   �h���Ë���j�)���Y����������������������������̋�U��f�} u�E (  �uh��h~��u�u�u������]�������������jh�(	�,���3ۋu9^��   j�ӿ��Y�]�9^��   h (  S��	VS���������}�;�uj��E�PhB	������3��   W����Y���u���N�u���t�>�8 u�  ��j�r���Y��;�tJ�^S�b���Y����t3�u�SV�+�����3�;�u�E�p�7�E�H�O�x�QQQQQ�X���W�O���Y�u��F���Y�u�E������   �F� ���Ëuj�����Y��������������������������������������������������������������������jh�(	�����j蒾��Y�e� �E�p��t�~�6����V����YY�����E������   �g����j�,���Y��������������������������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�������������������������������������̋�U��]�y����̋�U���V�u�M�������u�P�{�����e�F�P�Y�����Yu��P�^���Y��xu���M����   �	��	�F�����F��u�^8M�t�E��`p�������������������������������̋�U���V�u�M��T����E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p����������������������������������̋�U����E�����Az3�@]�3�]�������̋�U��QQ�} �u�ut�E�P�����M��E��M��H��EP�����E�M��������������������̋�U��j �u�u�u�������]������̋�V����tV覾��@PV�V�i�����^�������̋�U��j �u����YY]����̋�U��j �u�r���YY]����̋�U���SV�u�M��������3�;�u"����j^�0�V����}� t�E��`p���^[��9Mv�9M~�E�3���	9Ew	�v���j"��W8Mt�U3�9M��3Ƀ:-����ˋ��'����}�?-��u�-�s�} ~�N�E�����   � � F�3�8E��E��}�u����+�]h0�SV�l�������ut�N9Et�E�G�80t/�GHy���F-��d|�jd_�� F��
|�j
_�� F�� F�lo	_t�90uj�APQ��������}� t�E��`p�3������3�PPPPP�;�������������������������������������������������������������������������������������������̋�U���,�B	3ŉE��ESV�uW�}j[S�M�Q�M�Q�p�0�%�������u�������������m�E��t���u��3Ƀ}�-��+�3Ʌ���+��M�Q�NQP3��}�-��3Ʌ�����Q��������t� ��u�E�j P�u��V�u�������M�_^3�[�=�����������������������������������������������������̋�U��j �u�u�u�u�u�9�����]��������̋�U���$VW�u�M��E��  3��E�0   �����9}}�}�u;�u#�����j^�0�f����}� t�E�`p����  9}v؋E��� 9Ew	����j"�ȋ}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW�E�������t�}� � ��  �M�ap��  �;-u�-F�} �0����$�x�Fje��V����YY���U  �} ���ɀ����p��@ �;  %   �3��t�-F�]������$�x����0�F�O�����  �3���'3��u$�F0�O����� ���u�U���E��  ��F1����F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~L�W#U���M�#E���� �s���f��0����9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� � ���f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V������u�E�8 u���} �4����$�p���W����3�%�  #�+E�SY�x;�r	�F+����F-������ڋ��0;�|$��  ;�rSQRP����0�F�U�����;�u��|��drj jdRP�ݪ��0��U�F����;�u��|��
rj j
RP跪��0��U�F���]�0��F �}� t�E�`p�3�[_^������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �u�u�u�u�u�n�����]��������̋�U���SVW�u���w�ٍM�N�k�����u#�X���j^�0������}� t�E��`p����   �} v׀} t;uu3��?-���f�0 �?-��u�-�s�G��V�^芶��@PVS�O����0�������} ~QV�^�f���@PVS�+����E����   � � ������y&�߀} u9}|�}�}���u���Wj0S�������}� t�E��`p�3�_^[�����������������������������������������������������������������̋�U���,�B	3ŉE��EVW�}j^V�M�Q�M�Q�p�0�K�������u� ����0�������lS�]��u������0�������S���;�t3Ƀ}�-����+��u�M�Q�M��QP3��}�-���P��������t� ��u�E�j VS��������[�M�_3�^�e����������������������������������������������������̋�U��j �u�u�u�u������]�������̋�U���,�B	3ŉE��EV�uWj_W�M�Q�M�Q�p�0�6�������u������8�������   �M��t�S�]�3�K�}�-���<0���u��+ȍE�P�uQW��������t� �W�E�H;������|-;E}(��t
�G��u��G��u�E�j�u���u���������u�E�jP�u���u�u�y�����[�M�_3�^�$���������������������������������������������������������������̋�U��j �u�u�u�u�u������]��������̋�U��E��et_��EtZ��fu�u �u�u�u�u�z�����]Ã�at��At�u �u�u�u�u�u�X����0�u �u�u�u�u�u�O�����u �u�u�u�u�u膥����]����������������������������������̋�U��j �u�u�u�u�u�u������]��������̋�VW3��� B	�ܑ	�� B	����(r�_^��������̋�Vh   h   3�V��������t
VVVVV�y���^�����������j
���	���	3������j �ܑ	������	� �̋�U���u�5TB	� �	��]� �����̡PB	Ë�V�5TB	� �	����u�5x_	�ԑ	��V�5TB	��	��^�������������̋�U���u�u�5|_	�ԑ	��]� ������̡PB	���tP�5�_	�ԑ	�ЃPB	��TB	���tP��	�TB	��������������������jh�(	�h���h8���	�u�F\���f 3�G�~�~pƆ�   CƆK  C�Fh�E	j����Y�e� �vh��	�E������>   j�ŭ��Y�}��E�Fl��u��N	�Fl�vl����Y�E������   �����3�G�uj�_���Y�j�V���Y���������������������������������������������̋�VW��	�5PB	���8����Ћ���uNh  j�������YY��t:V�5PB	�5|_	�ԑ	�Ѕ�tj V�_���YY�Б	�N���	V����Y3�W��	_��^������������������������������̋�V蕤������uj�,���Y��^�������jh)	������u����   �F$��tP����Y�F,��tP����Y�F4��tP����Y�F<��tP����Y�F@��tP�u���Y�FD��tP�g���Y�FH��tP�Y���Y�F\=��tP�H���Yj����Y�e� �~h��tW��	��u���E	tW����Y�E������W   j�Ϋ��Y�E�   �~l��t#W����Y;=�N	t���M	t�? uW�a���Y�E������   V�����Y菾��� �uj�O���YËuj�C���Y���������������������������������������������������������������������������̋�U��=PB	�tK�} u'V�5TB	�5 �	�օ�t�5PB	�5TB	���ЉE^j �5PB	�5|_	�ԑ	���u襻���TB	���t	j P��	]�����������������������������%Б	�%�	��Wh8���	����u	蟷��3�_�V�5 �	h��W��ht�W�t_	��hd�W�x_	��hX�W�|_	�փ=t_	 �5�	��_	t�=x_	 t�=|_	 t��u$� �	�x_	��	�t_	r��5|_	��_	���	�TB	�����   �5x_	P�օ���   �}����5t_	�5ܑ	���5x_	�t_	���5|_	�x_	���5�_	�|_	�֣�_	�F�����tc�=ԑ	hR��5t_	���УPB	���tDh  j�������YY��t0V�5PB	�5|_	���Ѕ�tj V����YY�Б	�N��3�@��B���3�^_����������������������������������������������������������������������������������������������̋�U��V�uV�$�	���  ;5�_	v�����^]���������̋�U��M��_	��_	]�����̋�U��VW3��u�b�����Y��u'9�_	vV�$�	���  ;�_	v��������uʋ�_^]�����������������̋�U��VW3�j �u�u�\���������u'9�_	vV�$�	���  ;�_	v��������uË�_^]�������������������̋�U��VW3��u�u�k�����YY��u,9Et'9�_	vV�$�	���  ;�_	v��������u���_^]�������������������̋�U��VW3��u�u�u�N���������u,9Et'9�_	vV�$�	���  ;�_	v��������u���_^]��������������������̋�U��h����	��th��P� �	��t�u��]����������̋�U���u�����Y�u�(�	�������j葦��Y���j�^���Y��̋�V�������V�%���V����V萳��V����V菨��V������^������������̋�U��V������t�Ѓ�;ur�^]�������̋�U��V�u3����u���t�у�;ur�^]���������̋�U��M��u�U����    �����jX]á�_	��t�3�]������������̋�U��M��u�����    ����jX]á�_	��t�3�]������������̋�U��=<� th<�����Y��t
�u�<�Y����h@�h$��+���YY��uTVWh���a���� �� �Y��;�s���t�Ѓ�;�r�=��	 _^th��	�1���Y��tj jj ���	3�]��������������������������������������j h8)	�����j諤��Y�e� 3�@9�_	��   ��_	�E��_	�} ��   �5��	�5ԑ	�֋؉]Ѕ�th�5��	�֋��}ԉ]܉}؃��}�;�rK�ǫ��9t�;�r>�7�֋�贫������5��	�֋��5��	��9]�u9E�t�]܉]ЉE؋��}ԋ]���E�D��}�P�s�E� ��t�ЃE����E�T��}�X�s�E�� ��t�ЃE����E������    �} u)��_	   j�t���Y�u�'����} tj�^���Y�芶����������������������������������������������������������������������������������̋�U��j j �u�_�����]�����̋�U��j j�u�D�����]������jj j �/���������jjj ���������̋�U�������u�y���Yh�   �����������̋�U���LV�E�P�<�	j@j ^V�?���YY3�;�u����  ��   ���	�5T�	;�s6���H��f�@� 
�Hf�@ 
�@!
�H3�H/�5��	��@�P���   ;�r�SWf9M��  �E�;��  ����E�þ   �E�;�|��9T�	}k���	j@j ����YY��tQ�T�	 ��   �;�s1���H���` �`��`3 f�@� 
f�@ 

�@/ ���@΍P�;�r҃�9T�	|���T�	3���~r�E�� ���t\���tW�M��	��tM��uP�8�	��t=����������4���	�E�� ��E�� �Fh�  �FP�4�	����   �F�E�G�E�;�|�3ۋ���5��	����t���t�N��q�F���uj�X�
�C�������P�0�	�����tB��t>W�8�	��t3%�   �>��u�N@�	��u�Nh�  �FP�4�	��t,�F�
�N@�����C���h����5T�	�,�	3�_[^�Ã����������������������������������������������������������������������������������������������������������������������������������������������������̋�VW���	���t6��   ;�s!�p�~� tV�@�	���@   �N�;�r��7������' Y������	|�_^��������������������̃=��	 u�$���V�5T_	W3���u����   <=tGV�E���Y�t���u�jGW�������YY�=�_	��tˋ5T_	S�3V�����>=Y�Xt"jS����YY���t?VSP���������uG���> u��5T_	�����%T_	 �' ���	   3�Y[_^��5�_	�����%�_	 �����3�PPPPP�ӷ���������������������������������������������������������̋�U��E��_	]���̋�U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�v���Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#葰��Y��t��M�E�F��M��E���n���Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��������������������������������������������������������������������������������������������������������̋�U���S3�VW9��	u�����h  ��_	VS��`	�D�	�̄	�5�_	;�t�E�8u�u��U��E�PSS�}������E���=���?sJ�M���sB�����;�r6P������Y;�t)�U��E�P�WV�}��c����E���H��_	�5�_	3�����_^[�����������������������������������������������̋�U���SV�P�	��3�;�u3��wf93t��f90u���f90u�W�=L�	VVV+�V��@PSVV�E��׉E�;�t8P�4���Y�E�;�t*VV�u�P�u�SVV�ׅ�u�u��$���Y�u�S�H�	�E��	S�H�	3�_^[��������������������������������������̋�V��#	��$	W��;�s���t�Ѓ�;�r�_^���������̋�V��%	��&	W��;�s���t�Ѓ�;�r�_^����������j h   j �T�	3Ʌ����a	�����������5a	�X�	�%a	 �����̡a	�����h��d�5    �D$�l$�l$+�SVW�B	1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�����������������������̋���t�O�30�ڿ���O�G�30�ʿ�������������̋�U���S�]V�s35B	W��E� �E�   �{���t�N�38腿���N�F�38�u����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���K����E���x@G�E��؃��u΀}� t$����t�N�38�����N�V�3:�����E�_^[��]��E�    �ɋM�9csm�u)�=H�	 t hH�	螴������t�UjR�H�	���M�U�۵���E9XthB	W�Ӌ��{����E�M��H����t�N�38�l����N�V�3:�\����E��H��薽�������9S�O���hB	W���&���������������������������������������������������������������������������������������������������������̋�V9t�����   ;�r���   ^;�s9t3����������̋�U��V���������2  �N\�U��W9t�����   ;�r���   ;�s9t3���t�P��u3���   ��u�` 3�@��   ����   �MS�^`�N`�H����   j$Y�~\�d9 �����   |� �~d=�  �u	�Fd�   �~=�  �u	�Fd�   �n=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=� �u	�Fd�   �=� �u�Fd�   �vdj��Y�~d��` Q��Y�^`[���_^]����������������������������������������������������������������������������������̋�U��csm�9Eu�uP�k���YY]�3�]��������̋�U����B	�e� �e� SW�N�@��  ��;�t��t	�УB	�eV�E�P���	�u�3u��d�	3��Б	3��`�	3��E�P�\�	�E�3E�3�;�u�O�@����u��G  ����5B	�։5B	^_[���������������������������������������̋�U��} u� ����    �ķ�����]��uj �5a	�h�	]�������������f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U������������������������������������������������̋�U��E���#��	�<�	]�������j
���	�<�	3������U�������$�~$�   ��fD$f��f%�f-00f=��B  f���Y�f���-��X�f���\�f(���Y�fɁ�v ����?f(-��������fY��\��Y���\�fxf����\�fY�f\�f(5���Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-���Y fX5��fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f��\�fL$�D$����F����I �������������������������������������������������������������������������������������������������������������������̀zuf��\���������?�f�?f��^���٭^������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp��������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-����p��� ƅp���
��
�t���������������������������������������������������������������������������������������������������������������������������������������������ËT$��   ��f�T$�l$é   t�   ��0��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   贤��Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t�V���Z�萚��Z��,$Z��\������������L������   s��l���T������������D������   v��d������������������������������������������������������������������������������������������������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�C������E�f�}t�m�������������������������������U�������$�~$�   ��fD$f%0�f@�fW�f8���fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU��fV�f($������X��\��Y��Y��Y����X��^�f=��f-���\�fs�?��fs�?�Y�fp�Df5���Y��Y���fW��Y��Y��X��Y��X�fp���X��X��X�fD$�D$���-�  ��C�  �Y��\��Q�f��fs�fT=��fs���f%@����\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<����Y�f(���Y��Y��\��X��\��X�f-���\��X�f���^�f��f\ՠ����Y�%�   ���Y��Y΃��Y��Y��X�f���Y��X�f���X�fp���\��X�fV�fD$�D$����;  = 8  sjf�f(5��f�f( �f(%�fY���fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X�fD$�D$���-�;  ���O  �Y��\��Q�f��fT=��fp�DfT����f%@����\��Y��X��Y��\����Y��Y��\��\��X��\�f(��fp���\��X�fp���X��Y��X�fp���^�f( �f(- �f(�fY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f(���Y�fX�fp���Y��fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fV�fD$�D$����� = � ��   f~�fs� f~�����  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$�Y���fD$����fD$�D$���f0�f��f���X�fU�fV���fD$�D$���fD$fW��Xƺ�  �t���fD$fW�����f�����  �����  r�X�fV��Y�fD$�D$������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��3��M;�P�t
@��r�3�]Ë�T�]���������̋�U����  �B	3ŉE�SV�uWV������3�Y�����;��l  j�K���Y���  j�:���Y��u�=`_	��   ���   �6  h��h  �a	W臨��������   h  �Ba	VSf�Jc	�p�	��  ��uh��SV�O�������t3�PPPPP����V�*���@Y��<v*V�����E�`	��+�j��h��+�SP蘣������u�h���  VW�Py������u������VW�<y������u�h  h(�W�4������^SSSSS�y���j��0�	��;�tF���tA3��G�����f9Gt@=�  r�S�����P�����P�]�����YP�����PV�l�	�M�_^3�[�B����������������������������������������������������������������������������������������������������������������j�e���Y��tj�X���Y��u�=`_	uh�   ����h�   �����YY��������������̋�U��E3�;ͰB	tA��-r�H��wjX]ËʹB	]�D���jY;��#���]�������������������z����u�D	Ã�������z����u�D	Ã�����̋�U��V�����MQ��'���Y�������0^]��������̋�U���bz����ujX]������M�3�]��������̋�U��V�u��u
�o���jX�趤��� �3�^]���������̋�U���z����ujX]��`����M�3�]��������̋�U��V�u��u
����jX��3���� �3�^]���������̋�U��E�th	]���̋�U��Vj躁��Y�5th	�ԑ	�u���ܑ	j�th	�n���Y��^]��������������j �
���Y����5th	�ԑ	���̋�U���5th	�ԑ	��t�u��Y��t3�@]�3�]�����������W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y�������������������������������������������������������������������̋�U��} u	�%|h	 ]��u�ܑ	�0�	�|h	   ]�����������̋�U���(3��E��E�9|h	t�50�	�ԑ	�����M��   V;���  ��  ���  �  jZ+���   I��   ����   I��   ����   ItN��	�  �E�   �E����M��M�u�]���M��]�Q��]���Y����  �l���� "   ��  �E����M��M�u�]���M��]�Q��E�   �]���Y�  �E�   �E�����E����M�u��M�]���]���?  �U��E����W����E����ΉU��E����?����E����q�����tWItHIt9It ��t���  �E�����E�����E����M��u��u����E����c����E�   �������E���   �E�   �Eܸ��������������   �$�PN�E�����E�����E�����Eܰ���Eܨ��t����Eܠ��h����Eܘ��\����Eܔ���Eܐ���E܌��M��u�M����M�]���]�M��]�Q�E�   ��Y��u襟��� !   �E��^�Ð�M�M�M�M�M�M_M�M@M7M�M�MN����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��QQSV���  V�5lD	�O����EYY�M�ظ�  #�QQ�$f;�uU����YY��~-��~��u#�ESQQ�$j��}�����tVS�����EYY�f�ES������\$�E�$jj�A�}���]��E�Y�EY������DzVS辄���E�YY�"�� u��E�S���\$�E�$jj�w����^[�������������������������������������������������������̋�U���(  ��i	��i	��i	�|i	�5xi	�=ti	f��i	f��i	f�pi	f�li	f�%hi	f�-di	���i	�E ��i	�E��i	�E��i	��������h	  ��i	��h	��h		 ���h	   �B	�������B	�������̑	��h	j�v���Yj ���	h���|�	�=�h	 uj�R���Yh	 ��x�	P�t�	������������������������������������������������������������������̋�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H臆����t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�A����EPSj �u���	�M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��j �u�u�u�u�u�u�%�����]��������̋�U��j�u�u�u�u�u�u�������]��������̋�U����ESV3ۋ���C�u��t�]tS�'���Y����  �t�Etj����Y����x  ����   �E��   j�����EY�   #�tT=   t7=   t;�ub��M�����E	��{L�H��M�����{,��E	�2��M�����z��E	���M�����z��E	���E	��������   ���   �E��   3��t��W�}���������D��   ��E�PQQ�$�r���M��]�� �����������}�E���(��S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj蔇��Y�e���u��Et�E tj �y���Y���3���^��[��������������������������������������������������������������������������������������������������������������������������̋�U��}t~�}������ "   ]������ !   ]�����������̋�U��3���pD	;Mt
@��|�3�]Ë�tD	]���������̋�U��E� tj��t3�@]ètj��tjX]������]�������������̋�U��� 3���pD	;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���{���E�P�������uV��x��Y�E�^�Ë�tD	�h��  �u(�{���u�x���E �������������������������������������������̋�U��= Q	 u(�u�E���\$���\$�E�$�uj�ц����$]��i���h��  �u� !   �{���EYY]���������������������̋�U��QQ�= Q	 �E�E�]�u)�u�E����\$�E�\$�E�$�uj�[�����$������h��  �u� !   �z���E�YY�������������������������̋�S��QQ�����U�k�l$���   �B	3ŉE��s �CP�s��������u#�e��P�CP�CP�s�C �sP�E�P��{�����s��������= Q	 u+��t'�s �C���\$���\$�C�$�sP腅����$�P��v���$��  �s ��y���CYY�M�3�������]��[��������������������������������������������������̋�S��QQ�����U�k�l$���   �B	3ŉE��s(�C P�s��������u2�E��C����]����E�j �C P�CP�s�C(�sP�E�P��z�����s�������= Q	 u,��t(�s(�C ���\$�C�\$�C�$�sP�y�����$�P��u���$��  �s(�x���C YY�M�3��ڕ����]��[������������������������������������������������������̋�U��QQ�E�E�M�]��  �����  �f�E��E�������������̋�U���E��%�  -�  �]������̋�U���E�E�M��%�  �����PQQ�$�D�����]�����������̋�U��QQ�M�E�E�]������  �f�E��E������������̋�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]�f�M��  V��f#�^f;�uj���  f;�u�E�� u9Utj��3�]�������������������������̋�U���E������������Dz3��   �E3ɩ�  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$�������&Q���EQQ�$�ݏ���U�����  �����  �E�]������������������������������������������������̋�U��Q��}��E������̋�U��Q�}����E������̋�U��Q��}��E�M#M��f#E�f����E�m�E������������̋�U��QQ�M��t
�-�E	�]���t����-�E	�]�������t
�-�E	�]����t	�������؛�� t���]�������������������������̋�U��Q�=��	 t�]���e� �E����������jhX)	�T���3�9��	tV�E@tH9�E	t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�E	 �e��U�E�������e��U�~������������������������������̋�U��Q�=��	 t�]��e���U����������3�9��	t��j����?�����3�9��	t�j����?�I|��������̋�U��V3�95��	t"�j���M#M���E�����#��P�5g��Y��^]�������������̋�U���Qj���M��?�P�
g��Y]���������������������U���0���S�ٽ\�����= Q	 t�|����8����   [����ݕz������U���U���0���S�ٽ\����= Q	 t�D|����8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8�����{���   [�À�8�����=L_	 uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ��������������x�����s4����,ǅr���   ��������������p�����v���VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�6u����_^�E�����U���0���S�u�u�   ���ٽ\�����8�����lz������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�����������������������������������������������������������������������������������������������������������������������������������������������������������������a����tj�_{��Y��E	tjh  @j�)�����j�i��������������̋�U��M��E	�U#U��#�ʉ�E	]��������̋�U���   �B	3ŉE��}�ESVW�}��x�����   ��t��� h�   ��|�����Q�u�uP�4^��������ub��	��zuxVV�u�u��x����^������p�����tXFVP�f�����YY��tH��p�����t���S�u�u��x�����]��������tjV�/����3�YY;�u!9�t���tS袇��Y����M�_^3�[贌���ÍN�QSVP��`������u9�t���tS�n���Y3���WWWWW�b���}uH�5��	3�PP�u��u�֋؅�tjS謊��YY���tSP�u�u�օ�u��7�����' Y�p����} �f�����x��� j��x���P�E    P�u���	���<�����x�����c�������������������������������������������������������������������������������������������������������������̋�U��E�Dl	]���̋�U��QV�uV�Wr���E�FY��u�n���� 	   �N ����/  �@t�S���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,��v���� ;�t�v����@;�u�u�p��Y��uV��x��Y�F  W��   �F�>�H��N+�I�N;�~WP�u�a�����E��M�� �F����y�M���t���t�������������	��`B	�@ tjSSQ�m��#����t%�F�M��3�GW�EP�u�a�����E�9}�t	�N �����E%�   _[^��������������������������������������������������������������������������������������������A@t�y t$�Ix��������QP�}��YY���u	��������������̋�U��V����M�E�M�����>�t�} �^]���������̋�U��QSV�����R����G@� �E�t
� u�J�8����  �(�E� ��K�U����E�>�u�����8*u�ϰ?�:�����������8 u
������M��^[������������������������������̋�U��E� � �@�]����̋�U��E� ��A��Q�]�����̋�U��E� � f�@�]����̋�U���x  �B	3ŉE�S�]V�u3�W�u�}�������������������������������������������������������������.p����u+�����    迄�������� t
�������`p������
  �F@u^V��n��Y�`B	���t���t�ȃ����������	����A$u����t���t�ȃ��������	����@$��q���3�;��g����3ɉ��������������������������9
  G������9������&
  �B�<Xw���������3������j��Y������;���	  �$��t��������������������������������������������	  �� tJ��t6��t%HHt���u	  �������i	  �������]	  �������Q	  �������   �B	  �������6	  ��*u,���������[�������;��	  �������������	  ������k�
�ʍDЉ�������  ��������  ��*u&���������[�������;���  ��������  ������k�
�ʍDЉ������  ��ItU��htD��lt��w��  ������   �r  �?luG������   �������W  �������K  ������ �?  �<6u�4u�������� �  �������  <3u�2u�������������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������ ������P��P��^��Y��������Yt"�����������������G�������������������������������h  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@�������   ������������9������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  �������[���������  ;�u��E	������������ǅ����   �y  ��X��  HHty+��'���HH��  ��������  ������t0�C�Ph   ������P������P�ʀ������tǅ����   ��C�������ǅ����   �������������/  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ��E	������P�Y_��Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�3����������m�����:��������� tf������f���������ǅ����   ��  ������@ǅ����
   �������� �  ��  ��S����  u��gucǅ����   �W9�����~�������������   ~=��������]  V�rR��������Y��������t���������������
ǅ�����   ��5ԑ	���������C�������������P��������������������P������������WP�58B	���Ћ���������   t������ u������PW�5DB	����YY������gu��u������PW�5@B	����YY�?-u������   G������W�
���ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �p���������Qƅ����0������ǅ����   �L�����   �R������� t��������@t�C���C����C���@t��3҉�������@t��|��s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�d����0���������ڃ�9~������N뽍E�+�F������   ������������tb��t�΀90tW�������������0@�?If90t��;�u�+��������(;�u��E	�������������I�8 t@;�u�+����������������� �}  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+������������u'����~!������������� O�����������t��ߋ�����������������P�����������������Yt(������u��������ϰ0K�W����������t��ヽ���� ������tT��~P�������Pj�E�P������PK���U{������u ��������t�E�P�������e���Y��u�������������������������B���Y������ |.������t%��������������ϰ K�����������t��ヽ���� t�������x�������� Y���������������t������������3�������������� t
�������`p��������M�_^3�[��|���ÍI �l�jk_k�k�k�k-m��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��E�Hl	]���̋�U���(  �B	3ŉE�S�]W���tS�_[��Y������ jL������j P�(R����������������0�����������������������������������������������f������f������f������f������f������f��������������E�M������ǅ0���  �������I��������M�������M�������������̑	j �����	������P�|�	��u��u���tS�jZ��Y�M�_3�[�x�����������������������������������������������������������������������������̋�U��V�5Hl	�ԑ	�u���ܑ	�Hl	��^]�����������5Hl	�ԑ	���̋�Vj� �Vj�Oo����V�x�	P�t�	^���������̋�U���u�u�u�u�u�j��������̋�U���5Hl	�ԑ	��t]���u�u�u�u�u�}j��������������3�PPPPP� k���������3�VPPPPP��j��j� �Vj�n���� V�x�	P�t�	�����������̋�U��]�j����-�  t"��t��tHt3�ø  ø  ø  ø  �����������̋�VW��h  3��FWP�O��3��ȋ��~�~�~����~�����E	���F+ο  ��@Ou���  �   ��@Nu�_^�������������������������̋�U���  �B	3ŉE�SW������P�v���	�   ����   3�������@;�r�����ƅ���� ��t0���������;�w+�@P������j R�N�����C����u�j �v�������vPW������Pjj �a��3�S�v������WPW������PW�vS�b����DS�v������WPW������Ph   �vS�b����$3���E������t�L���������t�L ��������  ���  @;�r��R��  ǅ��������3�)�������������  ЍZ ��w
�L�Q ���w�L �Q����  A;�rƋM�_3�[��t��������������������������������������������������������������������������������������������������������jhx)	�hd����Y�����L	�Gpt�l t�wh��uj �j��Y���a���j��M��Y�e� �wh�u�;5J	t6��tV��	��u���E	tV��n��Y�J	�Gh�5J	�u�V��	�E������   뎋u�j�fa��Y�����������������������������������������̋�U���S3�S�M���[���Ll	���u�Ll	   ���	8]�tE�M��ap��<���u�Ll	   ���	�ۃ��u�E��@�Ll	   ��8]�t�E��`p���[��������������������������������̋�U��� �B	3ŉE�S�]V�uW�E�����3��};�u�������3��  �u�3�9� J	��   �E��0=�   r����  �t  ����  �h  ��P���	���V  �E�PW���	���7  h  �CVP�K��3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP��J���M��k�0�u���0J	�u��+�F��t)�>����E���J	D;�FG;�v�}���> uЋu��E����}��u�r�ǉ{�C   ����j�C�C��$J	Zf�1f�0����Ju���+��������L@;�v����~� �0����C��   �@Iu��C�A����C�S��s3��ȋ�����{����95Ll	�T�������M�_^3�[�=q�����������������������������������������������������������������������������������������������������������������������������̋�U���j �M���X���E�x t�}� �@t�M��ap��À}� t�E��`p�3������������������jh�)	�P`���M����U�����}��0c���_h�u�����E;C�W  h   ��@��Y�؅��F  ��   �wh���# S�u�J��YY�E�����   �u��vh��	��u�Fh=�E	tP��j��Y�^hS�=�	���Fp��   �L	��   j�]I��Y�e� �C�\l	�C�`l	�C�dl	3��E��}f�LCf�EPl	@��3��E�=  }�L��H	@��3��E�=   }��  ��I	@���5J	��	��u�J	=�E	tP�j��Y�J	S���E������   �0j�\��Y��%���u ���E	tS��i��Y�k���    ��e� �E��[��������������������������������������������������������������������������������������������������������̃=��	 uj���l��Y���	   3��������̋�U��SV�5�	W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�L	t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]�����������������������������������̋�U��W�}����   SV�5�	W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�L	t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]��������������������������������������̋�U��SV�u���   3�W;�to=8T	th���   ;�t^9uZ���   ;�t9uP�{g�����   �qa��YY���   ;�t9uP�Zg�����   �a��YY���   �Bg�����   �7g��YY���   ;�tD9u@���   -�   P�g�����   ��   +�P�g�����   +�P��f�����   ��f�������   = L	t9��   uP�^f�����   ��f��YY�~P�E   ��L	t�;�t9uP�f��Y9_�t�G;�t9uP�f��Y���Mu�V�vf��Y_^[]����������������������������������������������������������������������������������̋�U��W�}��t;�E��t4V�0;�t(W�8�`��Y��tV�a���> Yu���M	tV�gl��Y��^�3�_]��������������������jh�)	�Z���OP����L	�Fpt"�~l t�8P���pl��uj ��`��Y���RW���j�?D��Y�e� �5�N	��lV�b��YY�E��E������   �j��W��Y�u�������������������������������̋�U��UVW��t�}��u�Hf��j^�0��f�����3�E��u����+���@��tOu��u� �f��j"Y�����3�_^]�����������������������̋�U��E��u��e���    �f��jX]Ë�N	�3�]�����������̋�U��E��u�e���    �Gf��jX]Ë�N	�3�]�����������̋�U��E��u�ke���    �f��jX]Ë�N	�3�]�����������̋�U��S�]V��t4�} v4��t� W�}��t�E��t1��t,�e��j^�0�e�����K�} t���d��j^�0�e�����3�4�xO	�6�iE��@Y���u3��;Evj"X��6�uS�,f����_^[]������������������������������������̸�N	ø�N	ø�N	øxO	Ë�U���1h���M�]����̋�U���QQ���M�]����̋�U���eZ���M�]�����j,h�)	��W��3ۉ]ȉ]ԉ]�]܉]؉]�j�A��Y�]��B���E��E�P�M��Y;���   �E�P��I��Y;���   �E�P�T<��Y;���   ��>���Ẻm	����=�O	�=�O	hl��l:��Y���u�;�tt8tp� m	;�t!PV�{D��YY���A  � m	;�tP�5b��YV��C��@P�8��YY� m	;��  VV��C��Y@P�5 m	�d����;���   SSSSS��Y��� m	;�tP��a��Y� m	hpl	���	;���   3�A�m	�pl	k�<�E�f9�l	t��l	k�<E�f9
m	t�m	;�t�M�+�l	k�<�E���]܉]؍E�PSj?�E��0Whtl	S�ű=L�	�ׅ�t9]�u
�E�� �X?��E�� ��E�PSj?�E��pj�h�l	S�u��ׅ�t9]�u�E��@�X?��E��@��E�   �}��RX���8�}���e���8�}��O���8�E������Y   9]���   jVj@�}��7��9��������������>-u�E�   FV�a��Yi�  �E�<+t<0|<9F��3ۋu�j�S��YÀ>:u8FV��`��Yk�<E��<9F�<0}��>:uFV�`��YE��<9F�<0}�9]�t�]���E�;�tjVj@�w�Y9������t
�����G��u��YW���0�u���d���0�Q������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����e� �}SVW�}������   %  �yH���@�E�u��jd�[����u��l  ���  ����t�������T	��������T	�E��+  ��_���  ��jd_Fj�E��Ù���U��}[+ЉU��G��������E���i�m  ��%�������Ek�+�E;U�t����}��   �}� u��jd�[����u��l  ���  ����t�E���T	�	�E���T	;�~D���?%  �yH���@u��jd�[����u��l  ���  ����t	�4��T	��4��T	uk�<M k�<M$i��  M(�}u�5�O	��O	�=�O	_^[�ÍE�P�5�O	��O	�<7��Y��uD�E�i��  �O	y��O	 \&��O	�� \&9�O	|)�O	��O	�=�O	�3�PPPPP�2U�������������������������������������������������������������������������������������������������������������������������������̋�U���V�E�3�P�u���C��Y����  9u��X  �WS3�C;�O	u;�O	�  95m	��   �m	�m	P�m	P�m	Pf95m	u�m	VP�m	PRS��m	PVVRV�
m	S�������l	��l	��$P��l	P��l	Pf95�l	u��l	VP��l	P�wS���l	PVV�wV��l	V������$�TjXjY�E�   �]���k}jX���E�
   �E�   VVVVVQRSSjY�K����E�VVVVV�u��wSVjY�3�����H��O	��O	�W;�};�|";�;�~;�}��[^��;�|�;��;�~;�}3���Gk�<Gk�<i��  ;�u3�;�O	���3�;�O	�����VVVVV��R������������������������������������������������������������������������������������������������������������������������jh�)	�dO��3�95$m	u*j�9��Y�u�95$m	u�;����$m	�E������   ��K���j�L��Y��������������������jh*	�O��j�8��Y�e� ������E������   �K���j�lL��Y���������������jh8*	�N��j�q8��Y�e� �}������E��E������	   �E��XK���j�L��Y����������������̋�U��UV�uW��H�F��w�� �
�y�B��w�� ��t;�t�_+�^]��������������̋�U���S�u�M��VF���]��u#�@Z���    ��Z��8]�t�E��`p������V�u��u$�Z���    �Z���}� t�E��`p������R�E��x uVS�]8��YY�1+�W�3�M�QP�9������M�QP��8����F��t;�t�+���_�}� t�M��ap�^[�������������������������������������������������̋�U��3�9�o	u'9Eu�WY���    ��Y������]�9Et�]�7��P�u�u�kI����]�����������������̋�U����u�M��E���E�M����   �A% �  �}� t�M��ap����������������̋�U��j �u�6��YY]����̋�U��h  �u�E��YY]�����̋�U��h  �u�yE��YY]�����̋�U��j�u�aE��YY]����̋�U��j�u�JE��YY]����̋�U��j�u�3E��YY]����̋�U��j�u�E��YY]����̋�U��j�u�E��YY]����̋�U��j�u��D��YY]����̋�U��h�   �u��D��YY]�����̋�U��h�   �u�D��YY]�����̋�U��j�u�D��YY]����̋�U��j�u�D��YY]����̋�U��j�u�sD��YY]����̋�U��j�u�\D��YY]����̋�U��h  �u�BD��YY]�����̋�U��h  �u�'D��YY]�����̋�U��hW  �u�D��YY]�����̋�U��hW  �u��C��YY]�����̋�U��h  �u��C��YY]�����̋�U��h  �u�C��YY]�����̋�U��j �u�C��YY]����̋�U��j �u�C��YY]����̋�U�츀   f9E���]�����̋�U��h  �u�YC��YY��u	f�}_t]�3�@]���������̋�U��h  �u�*C��YY��u	f�}_t]�3�@]���������̋�U��h  �u��B��YY��u	f�}_t]�3�@]���������̋�U��h  �u��B��YY��u	f�}_t]�3�@]������������������������Q�L$+ȃ����Y�{/��Q�L$+ȃ����Y�e/������������̋�U����e� V�u��u�fU��j^�0�V�����  j$h�   V��1���E����tӋ�@�M��E���|��@W��s�U��j^�0뼃�|
���&A�w�SWj h�3�PQ��0���HF��+  ���  ���y�jd�}��M�؋Ǚ_��j�h����+؋E��������D��A��ڙRP��.��+��j ��Q SRP��.���}��U�}� M|��sG�E��ǀ3��U� �ȁ�  ��EyI���Aujd�Y����u�El  ���  ����uA��U� �2�E�ȁ�  �yI���Au
jd�Y����u�El  ���  ����u�E�   �Ej S�u�FW��/��j��F�h����RP�*.���U�}� ��T	u��T	�F3�A9B}��A9�|���Q I�N+�j �F�ES�p�0�/��j��Y���3�Sh  �u�W�V�o/��j��F�h����RP�-��S�U�j<�u�W�L/���Fk�<+��>_�^ 3�[^�����������������������������������������������������������������������������������������������������������������������������������������������̋�U��V�:������t�uV�I�����Y��Y#�^]������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� ������������������������������������������������������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� �������������������������������������������̋�U��Q�e� V�u��u�P��j^�0�VQ�����  Sj$h�   V�-���]����u�P��j^�0�(Q������@W��}�hP��j^�0����   ���W�������iҀ�y�ʍ�F   ��3�;�|+�B;�|+ȸ ��B;�|B+���E�   ���V���Q ����T	�Fi�����ȃ}� u��T	�F3�B9G}��B9�|��]J�V+���Q �F����j_j<�f  ��������  �V���_�Fi�����ȋ����_�Fk�<+ȉ3�[^���������������������������������������������������������������������������������̋�V�$������u�%O���    3�^Ã~D uj$��#��Y�FD��t܋FD^�������������̋�U��V��6������t�uV�E�����Y��Y#�^]������������������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� �������������������������̋�VW3��Pm	�<��O	u���O	�8h�  �0���4�	��tF��$|�3�@_^Ã$��O	 3��������������������̋�S�@�	V��O	W�>��t�~tW��W�xL���& Y�����P	|ܾ�O	_���t	�~uP�Ӄ����P	|�^[���������������������̋�U��E�4��O	���	]�������t$j ���	h�   �Z-��Y�������jhX*	��@��3�G�}�3�9a	u�E��j�M-��h�   � -��YY�u�4��O	9t���mj�!��Y��;�u��L���    3��Pj
�T*��Y�]�9u+h�  W�4�	��uW�oK��Y�L���    �]���>�W�TK��Y�E������	   �E��=���j
��=��Y������������������������������������������������̋�U��EV�4��O	�> uP�"��Y��uj�.F��Y�6���	^]������������̋��  Ë�U��E��E�A3��A�A�A]� ������̋�V��~ t��F� �v�F�VY�F�F��u�^����������̋o	���u3�À�0|��9��/A�o	�3�� ��t݀�A|*��P%���A�D¿�o	���@uۊA�o	��@t���������������������������̋o	SV� @  W3��9_u	A��o	�<A|<Z��   <$�1  2�A�o	���B��  ��  ����  ��$�T  �yPuAA�o	���J�n  �� �[  ��FtHH���L|y��M~��O�I  ��QufA�o	�\������A� �  A�o	�t��    �����������  ������   ��t
��������#�ȃ�tE��t#��t
���  �  ��t��?����<�������4��t�濁΀   �%��������   ���t�������@������������ �P  HHt*HHtHHu���������   �3  ��������   �"  ��t��������   �  #��  ��/�O�����5��   ��A�=����������� �  �y  ���  ��  A�o	�<0|<9���Dѣo	�<H��   �  ���  �9  ���  I�.  �� �  �#  ��C�  H��   H��   �������A�o	��<0��   <5��   �� �  ��0�   ��t
����������������t��������   ���������   �t��    ����������� t=HHtHH�1�����t��?����r�������j��t�濁΀   �[��������   �M��t�������@�>��������43Ʉ�������  �  �������� �  ��������� �  ��� |  A�o	�U  �<0�,  <8�$  ��A��Ё�����o	���y����$�}�� �  ��t��������   ���������t�������@��   ��������   ��   � �  ��t��������   ���������t�濁΀   �   ��������   �   � �  ��t��������   ���������t��?����w�������o��������e�������� `  �W��������    �I�������� h  �;�������� p  �-�������� x  �<9uA�o	���  �3Ʉ�������  ��_^[�W���צ� ��.�<�J�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̡o	�Ѓ���̡o	���Ѓ����̡o	���Ѓ����̡o	���Ѓ����̡o	���Ѓ����̡o	���Ѓ����̡o	��`3�<`��������̡o	���Ѓ����̡o	���Ѓ����̡o	��	�Ѓ����̡o	%   ��̡o	%    ��̡o	% @  ��̡o	���Ѓ����̡o	%   ��̡o	���Ѓ����̋�U��o	�Ш�E����u��]�������̋�U��VW�}������} ��tW�Y�d��uj_�FS;�sE�   ;�w8jh  ��n	��;����t�  �3���t�N��t���F+߉F�^�	3��+ǉF�F�N�D[_^]� ���������������������������������̋��  �@ �`� ������̋�U����M���I�H]� ������3��y�����3�9������AË��H   ��̋A�������3�9t
�A   t@����̃9 t�I   ����3�9t
�A   t@����́I   ��̋A������̋A������́I   ��̋A������́I    ��̋A������́I @  ��̋A������́I �  ��̋	��u3�Ë� ��̋	��u2�Ë�`��̋�U��	��u�E]� �]�`�����̋�U����xt�M�Q��~�P]� ������̋�U����M���I�H]� ������3��9	����̋���Ë�� ����̋�U����M� ���H]� �����3�@ÊAË�U��E;Es�I�@]� ����̋�U����M� ����t�Q��t��u3ɉH]� ���������̋A��t� ��t����"3������̋A��t� ��t����b2������̋�U��A��t� ��t���]�b�E]� �������̋�U��U���PJ��҃����� ���P]� ��������̋AÃy����$ ���̋�U��3�A�ho	u]	ho	���3ң,o	�0o	�4o	�8o	�<o	�@o	   �Do	�Ho	   �Lo	�Po	�To	   �Xo	�E��w
k�,o	]øPo	]���������������������������������̋�U����M�H��H�M� ���H]� �������̋�V��~ }�N�SW�~��؋����_�^[�F^����������̋�V��N��P��u	�N�^�`^�������̋�U��V�u��N�u��P;Es�u�N�P�R^]� �����������3�8t@A�9 u����̋�V���t+Ȋ�@Nu�^�����̋�U��} u3�]Ê��t:uAB�Mu���
+�]����������̋�U��U�����H,�	��o	�o	�U��tV�u�5o	�o	^��%o	 �%o	 ��n	�M�o	�M��n	�o	�o	 ]� ��������������������������̋�U���3ɸ  ��!E�!E�Q�E�PhR��E�P�u�M��M��aA���E�����������������̋�U����e� �e� �  ��!E�!E�j�E�PhR��E�P�u�A���E�����������������̋�U���u��n	�u��5��]�����̋�U��EV�uW�}+�;�~����t�E��+ǋ�S��AJu�[�7_^]�������������̋�U��} V��t0j j��n	�`5����t�u���J���3��������$�F��& �F �f� ����^]� �������������������̋�U��V��M�f� ����t	��t3�����& �F��uQ�~9��Y���u�F��^]� ����������������̋�U��S�ًV�uW��t<��u���xVW��n	�4������t&��}���u�����T>�RV�P�  ���t� _��^[]� ����������������������̋�U��VW�}���t.j j��n	�+4����t��H�� ���H�x�3����u�F_^]� �����������������̋�U��V��& �F �f� ���} t&j j��n	��3����t�u������3����u�F��^]� ������������������̋�U��EV��f� ���F��uP�8��Y���u	�F��& ��^]� ������������̋�U��V��>	t6W�}�? t,j j��n	�'3����t���O�H�3���t���D�_��^]� �����������������̋�U��E��	w1����t;��L���E��I�H� �E�`� ���  �@��Mj�,���E]� ������������������̋�U��VW�}��� 	��t1�} t+j W��n	�d2���F�~��t��t�M+Ȋ�@Ou���f �f _��^]� ��������������������̋AËA��t�I�D��2�����̋�U���q�q�u�u�:����]� ������̋�U��yujh 	�u�u�|:������E]� ���������̋�U��o	�8@�uu�M�o	�'���
�u�d��YY�E]������������̋�U���u����EY]����̋�U��V��~-�> �Et��t��t��tP��5��YP���-���P������^]� ���������������̋�U��SV��3�9t�f� ���F��_W�};�tR�E;�tK+�tAHS��n	tj��0��;�t%�u��W�� ���j�0��;�t�� ���H�3��;�u
�F��F_^[]� �������������������������������̋�U��3�V��F�f� ���8Etj�EP�'����^]� ����������̋�U��E3�V��V�f� ���;�t3�8tA8u�;�v	QP���>'����^]� ��������������̋�U��V�u3�W���W�g� ����;���   8��   �E��:EtK<_t<<$t8<<t4<>t0<-t,<a|<z~$<A|<Z~<0|<9~<�r<�v�o	   t;BA����8 u�R�u���&������t@�:Mt�' �G�� u
�G��G��_^]� ����������������������������������������������̋�U���$�B	3ŉE�S3�V��W�F�f� ���}���E�j j
�uO�u�y����0�E]���UuލE�+�PW����%���M�_��^3�[�9:���� ��������������������������̋�U���(�B	3ŉE��EV��3ɈN�f� ��W�}���M��M�;�|9Ms�U����E��؉US�3�Qj
P�uO������0�E��M��ȉ]�u�[8M�tO�-�E�+�PW���(%���M�_��3�^�9���� �������������������������������������̋�U��V�u�u��A�ΉF�<����^]� ��������̋�U��V��~.�E���u�@P���	����> u
��@�F�Q����)����^]� ���������������̋�U��W���RV�u��tI�? uV�'���<�F��t<t��P����&j j��n	��,����t
V�������3�P���a)��^��_]� ������������������������̋�U��3�V��F�f� ���8Etj�EP��#����^]� ����������̋�U��E3�V��V�f� ���3�8tA8u�QP���#����^]� ������������̋�U��QQ�o	� ����   ����A�o	��w�U��e� �� ��jYщU��o	������tK����� t0+�t)+�t!+�t+�t��t+�u*j�j�j�j�	j�Q�j�����P�M�����E�M���M��H�ËE�`� ���  �@�ËMj�o%���E���������������������������������������������������̋�U��o	� ��t,<At�E�`� ���  �@]ËM�o	h$ 	����
�Mj��$���E]������������������̋�U��V�u�u��A�ΉF������^]� ��������̋�U��V�u�u��A�ΉF��0����^]� ��������̋�U��V��~=S�]��t4�> uS� *���'j j��n	�O*����t� ���X�3�P����&��[��^]� �������������������̋�U��W���OSV�u3�;�tB8t>9uV�r���2Sj��n	��)��;�t3�8tB82u�RV�������3�P���T&��^[��_]� ������������������������̋�U���S3�V�u�^�f� ���E�   �8^��   W�o	� <@��   <Z��   9]�t�]��	j,���#4���=o	�:���   ����0��	w!��n	P�E�GP�=o	���P���C���Y�e�  ���E�P�E�P�]��	���o	+�YY��~��n	�9	t	�E�P����E�P������9=o	u�f� ���F�8^�8����	j���L��_��^[������������������������������������������������������������������̋�U��QQ�E�V�u��@h, 	�ΉF�`'���E�P��4��YP���V��j}����2���o	�8@u�o	��^����������������������̋�U��QQ�u�M��u�u�$�����j	���E����������̋�U��QQ�u�M��u�u�!�����=	���E����������̋�U��QQ�u�M��u�u������	���E����������̋�U��V�u�u��A�ΉF�%2����^]� ��������̋�U��V�u�u��A�ΉF�J&����^]� ��������̋�U��o	��S3ۀ9QuA�4 	�o	���u�Mj�� ���E�	  <0|L<9H���/�AR�o	P��t�M��$��P�E�SP�!������M��z$����M��@�A���   VW3�3��)��tI<A|2<P.������A�����A���o	�<@uӊA�o	<@t"�E�`� ���  �@�b�Mj�$ ���E�S�} WVt��t
�M���#����M���#���$��t�M���#��P�E�SP�� ������M��#����M��@�A��_^[����������������������������������������������������������������������������������̋�U����o	� �e� �e�  ������   ����Ѓ�w|�$�w�h| 	�ht 	�hl 	�hd 	�M�����o	� �o	��1tHHtHHtHHu$�E�P�E�PhX 	�M����������M��U���U��M��E��P�ËE�`� ���  �@�ËMj����E�Ð�������������������������������������������������������������������������̋�U��o	� ����X��   HH��   �E�P�1��Y�M���uh�o	� ��t]<@tS<Zt�E�`� ���  �@�áo	�o	���Ш�� 	u�� 	P�E�P�M�������M��@�A�����o	�E�U���H�áo	�o	���Ш�� 	u�� 	P��o	h� 	�M�����E���������������������������������������������������������̋�U��o	� ����tL<Zu�o	�U��E3Ɂ�  ����P�ÍE�P�s#��YP�E�Ph� 	�M��������}��j)�u�M��!j)�u�E�jPh� 	�M����������,��������E�����������������������������������̋�U���$�e�  ��S3�3��o	�o	���V����AW�� ���a  N�*  N�  :��  �o	�R:���   9]t�E�`� ���@�L  �o	�������t�Ѓ�vA�e� ����e�� ��j�E�P�M��E�,�]����SV�M����P�E�P�M��_����@��E��M�j>�M�E��,���o	�:$�E�M��E�M�u�o	��M�j^�M�E��V,���E�E�E��E��o	8t�o	�
j�M�� ���M��E�U�� @  ��H�v�Mj�4���E�g�E� \��K9]������E�e� ���!}�� j�E�P�M��E�>�]��:���9]u�M��8&�\�t�����E�o	�X!x�_^[�������������������������������������������������������������������������������������������������������������������̋�U��o	��8S3�8�B  �w���E�;�}�]�9]�u�E�j]P�E��M��  �e�  ��VW�}�   �]��wtfh$��M�����W�E��M���tS�o	8tJ�E�SP���YYP�E�Pj[�M�������R���E��E�E�j]�M�E��|*���E�P�M������}�~�9tn�wt�E�P�E�P�������M��@�MW�E�Pj(�M��8������ ���E��E��E�j)�M��E��*���E��E�E��E�E�P�M��^���E�E��E�E�E�P�E�P�����E�U�YY�M��_��H^�   �E9t`P�E�Pj(�M�������u ���E؉E�E�h� 	�M�E������E�E��E�j�M��E��X����E��E��E�j]�M��E��p)���E��$�E�j]P�EЍM�jPj[�T�����(�����m���P�u�1���EYY[������������������������������������������������������������������������������������������������������������������������������̋�U����E�j P���YYP�E�Pj`�M�������N���j'�u�M������E����������������̋�U��j�u�q���EYY]�����̋�U��j �u�V���EYY]�����̋�U��j �u�;���EYY]�����̋�U��E��� SV�u3ۉ�@C�F:��4  �o	�9 �  �E�P�E����E�Y�E��E�j �M��E���'��V�E�P�M��{������@�F:���   �o	�8@��   h, 	�o�o	� ��tp<@tl�E�P�u)��YP�E�Pj`�M��k�����%����E��E��E�j'�M��E��O'���E�P�������o	�8@u@�o	8^6�8@th� 	���p��8^~�8^�o	�8 uS�������j}����&���o	�8@u,�o	�$:� V�E�PS�M������������E���E�F��^[����������������������������������������������������������������������������������������̋�U����u�M������o	� �o	<@u|�o	� �o	<_uk�o	�E�j P�3���E�j P�(���o	�����t��@t@�o	���u�8 u�MHj�o	����E�ËM�@�o	�E��M��H�ËE�`� ���  �@���������������������������������������������̋�U��QQ�o	� ��u�Mj����/j <?u�o	�E�P�g��Pj-�u��	�����
�u�O��YY�E���������������������̋�U����   �B	3ŉE��o	S��o	V�uW����D�#  �u  �� �   ��0��   O��   Ou@�E�P�>&����x���P�2&���}�YY��   ��|�����   jd�E�P�M������u�f� ���& �F�6  �E��E�<-u�E��E��E�.��E�.��x���PVje��`���P�E�P��@����|������]������������  �o	�8@u�o	h� 	���M�����  ��8���P�N��YPVh����p����)����V�_%���  �o	j�������  ��E�x  �0�����J��   ��Qt;��R����j ��x���j P�����E�P�%����x������|������F�0  �E�P��$���o	 @  Yt*j�E�P�M������E�P�]��P�o	YY��tP�����E�P��x����M�P��Du'h� 	�S����������h� 	V��x����&	���   h4 	��j{�M�������H|%��J ��P���P�!��YP�M��!���j,�M��"����Ft,Ot	OtFOt#OuV��h���P�$��YP�M������j,�M��"����X���P��#��YP�M������j,�M��l"����H���P��#��YP�M�����j}V�M��q����V���Y�M�_��^3�[�#�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��o	3Ƀ�8��   9Mt7�8Xu2@�o	�E9u�Mh� 	�x����   Ph	�u�P���   �8Yu�u@�u�o	�y���YY�uV�u�E�VP�����FYY^� @  t$�E�P�E�Ph 	�M������������U��M���    t�E�P�E�Ph� 	�ӋM��U��E��H���uj�u�G�����E����������������������������������������������������������̋�U���u�u����EYY]�����̋�U���|�B	3ŉE�S3�V�u�^�f� ����o	�E�   8^��  W�  ���o	�:���  ��@��  9]�t�]��j,�������o	��ʃ�0��	w@�o	Q� o	�E�P�H����M  !}�E��]��Xu@�o	h� 	�M��!���  ��$u@8t�o	�E�P�5����   ��?��   �E�P�� ���o	 @  Ytgj�E�P�M�����E�P�>��P�o	YY;�tP됍E�P�E�Ph� 	�M��?����������E��E؋E�h� 	�M؉E��3���E؉E�E��]�E�P�E�Ph� 	�M���������z����E��EЋE�h� 	�MЉE������EЉE�E��!}čE�P�E�P�]��?���YY��@�M�E�o	+E���~� o	�9	t	�E�P�b����E�P������8^�J���_�M���^�o	3�[����������������������������������������������������������������������������������������������������������������������������������������̋�U���   �o	�S3۹  ��!M�!M�V3�@�]��]�o	��A��  �g  ;��]  ��/�J  ��1~[��9�<  �@��4�P��M�����9]�t(�E�P�E�Ph��M��Z�����������E؉E��E܉E��M��E��M��H^[��!M�]�8]t|��x���P����YP�E�Pj<�M������������E�P�M������M�;�t��P<>u
j �M����j>�M�����E;�t� �o	8u�M��E��M��x���@�o	S����p���SP������@���M��E��5o	;�t+�~�1u%�E�P�E�Pj~�M��/����������M��E�M��E�9]������E�P�M��b��������H�o	�Mj����E�������B��  ��  ��Z��  ��_��  �@�o	��O��   ��D��  ��9kt@;�t���/��  ��6~��8��  �@��4����M������@��4����*����@��4����M������M�� �  �U��E��A�����?t9��@�$  ��B�  ��C�  jhL��E�P������M����   ��@�o	;��������0��  Sh	�ǃ�T��  ��S��  ��P��  I�����I��  �@��4����M��F����o	� :�uj�u�M�������������0�m  ���d  �4�X��M������o	� �o	��0��   ��1t��΃��B  �o	�2����E��E�E��E�E�P�M��q���j,�E�P�E�P���Y���&���P�M��Q���j,�E�P�E�P�d��Y������P�M��1���j,�E�P�E�P�D��Y�������P�M�����j)�E�P�E�SP���YY�������P�M������j'�u�M����������E�SP�{����E�YY�E�E�j �M�E��a���E�E��E�E�E�P�M������M��O�@��4����M������S�E�SP�E����@���M��E�;�t�   t�E�`� ���@�������M��E�P�u�����������U|҃�V��   ��W~ă�Y��   ��_u��@�o	��A|���D~
��F~��J��@��4�(������@��4�(��M�������o	�8?u%�E�P�����YP�M�������o	�8@u�o	��E�P�{���YP�M�����h	�M�����M�E��M��&����@��4��������@��4��������3�F�@��4�4��M�����;������9]�������M�   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��o	��   �8?�+  �x$�!  �M���M����X����S� o	V�5�n	�M���n	�M�W�=�n	��n	����X����o	� o	�8?�E� u@�o	�E�P�E�jP�����j�E�jP�# ����@���E��M��u�o	�}� uf�E�P���YP�E�Pj<�M�������C����E�P�M�������M��t��P<>u
j �M��]��j>�M��S���} t�o	�8 t�o	�E�M�=�n	_�5�n	��M�^� o	�H[�ËE�`� ���  �@��������������������������������������������������������������������������������������̋�U���8�B	3ŉE�S�o	���V�u��0�uȃ�	w��n	PCV�o	��������  �e� W�  ��!}��?uJ�E�j P����YY��@�E�o	�M�@�o	��@�W  H3ɣo	8��AQ�M�������;  �L	�����E�   ���t:uAF�M�u��	�+�u���o	�0�<	j�ˋ�[���t	:uAFKu��	�+���   �o	���E�P����o	 @  Yt2j�E�P�M������E�P���P�o	YY�M��tP�����   �M�h8	������E�P�E�PV�M��|�����������EԉE܋E�h� 	�M܉E��p���E�P�M��l����?�} t�o	�8@u�M�3�#��o	�E�M��j@ho	�M������@�M�E�} _t��n	�9	t	�E�P������M�Eȉ�M�H�M�^3�[�n����������������������������������������������������������������������������������������������������������������������������������������̋�U���SV�uW3�S�E�j�^�� ��!~P��M������@���F:�u?�o	� :�t4<@t;V�E�Phd	�E�P�E�P���Y����������f������@�F�o	� <@u�o	�N:�t!~�F��?9uj���M����0V�E�Phd	�E�Pj�M��x �����u������������@�F_��^[���������������������������������������������������������̋�U���u�����EY]����̋�U��o	�� VW����3���G#�t�   t3��o	� �e� �  ��!u��o	�� ��   ��Tt^HtTHtJHtHt
Hu\h�	�Mh�	�F�E�P�����YP�E�Ph�	�M������������E��E��E�E��h�	�h�	�h|	�M�������e� !u��t�E��E��E��E�E�P�����Y�E�P�M��Y����M��E��M�H��M�o	hi	�����E_^���������������������������������������������������������������������̋�U��o	�8?u'@�8$uj�u�#��YY�"j j �u�o	�|���j j�u�������E]������������������̋�U���j �+�����P�M��X����o	�8 tP�@�o	����0t1HHt��uA�E�`� ���  �@�ÍE�P����YP�M��+����h� 	�M�����
j�M�����h�	�M������M��E��M��H����������������������������������������̋�U���XSVW3��  ��!u�}��^
���M��99t�A   �E�   u�}����  u�E�`� ���@�8�_  ����  uQj�u�������E�A  ����  u��E��I�'  �]��e� �  �   �   �M  3��]�!}�}�   ���E�����t%   �#���t��%   ;��  �}� ��t%   �#���t��%   =   ��  =   ��  �� @  t_�o	��������t7���Шt.�E�P����YP�E�Pj �M��)�����������E��E��E��E���E�P�b���YP�M������   �U��Å�t%   �#����,  9}��#  �E�j P�����YY�M�E�P�E�Pj{�E�P��������p���P�M������E�P������   Y�5o	u>�E�P�E�Pj,�M��}������7����E��E��E�h�	�M��E�� ���E�P�M�����h�	�M�� ���E�P�i����o	Y���������/  ���������  ���  �E�P�E�Pj �M�������������E��E��E�j �M��E������E��E��E��EčE�P�M��"����M��EĉM��E���  !u�!u�!u�!u�!u�3��}��}��}��}؉}Ћ�;�t%   �#�;���   ;�tw��%   =   u>�E�jP�v����EȉE��ẺEčE�jP�_����EȉE��ẺE��E�jP�H������;�t'��%   =   u�E�jP�&���YY�EȉE��ẺE�E�jP�����EȉE؋E�YY�E�3�9}�tF�}� t��%   =   t2�o	��`<`�E�Pt����Y��@�MЉE������YP�M�����o	��������t/���Шt&�E�P�E�P�E�P����Y���-�����M��@�E���E�P����YP�M��-���E�8 tA�}� t0�o	   u$P�E�Pj �M��#�����������E�P�M��k������@�M��E�!u�3��}�9}�tE�E�WP�_���YYP�E�Ph�	�M������������E�P�M�� ����o	   tA�M���  3�Wj��n	�����;�t�8�@ �`� �����E�WP�����YY��@�MȉE̋u��Å�t%   �%   ���  ����   ��%   =   uz�E�P�E�Ph�	�M��o�����������E�E��E�j,�M��E��	���E��E�EĉE�E�P�M��V����E�E��E�j,�M��E������E��E��E��EčE�P�M��(����.��tN��%   =   u@�E�P�E�Ph�	�M���������^����E��E��E�j,�M��E�����E�P�M�������h�	�M������E؉E��E�h�	�M��E������E�P�M������E�P�����YP�E�Pj(�M��.�����������E��E��E�j)�M��E�����E�P�M��`�����t��%   =   t�E�P�M��B����o	���Ш�E�Pt� ���YP�M��!��������YP�M������o	���Ш��  ����  �E��Mȉ�E�G�ẺM��E��  �u�M�������E�� |  ����   ��#с� h  u�E�P�u����YY�@�������   ��#с� p  tم�u|��#с� `  uOP�E�P�+����E�YY�E��E�j{�M��E�� ���E��E��E��EčE�P�M��B���h�	�u�M������������u��#�;�u�E�P�u�6����i�����t��#�-   ���% `  ���@���   ��t%   �#ƅ�t$�E��Ӂ�   +����B�����t
h�	�   �}� ��t	#�-   �% `  ���@����t%   �#ƅ�t%�E��Ӂ�   ��   ���B�����thX	�Q�}� ��t	#�-   �% `  ���@����t%   �#ƅ�t-�E��Ӂ�   ��   ���B�����th	�M�������}� u��#�= x  ������}� t��#�-   ���% `  ���@����t%   �#ƅ�tX�M���%   3�=   ����Ʌ�u�M�3�=   ����Ʌ�t'�E�P�E�Ph�	�M��d�����������M��E��R����E�P�E�P�O���YY��M��@�9����M�   3Ҿ   ��9U�t#�+��% `  ���@;��s  �o	��	�Ш�M  ��9U�t#�+��% `  ���@;�tG9U�t��%   -   ���@�3�@;�t(�E�P�E�Ph	�M��������"����M��E��M��E�U���t��%   =   ��   ��t��#�+����% `  ���@����t%   �%   ����   �Å�t#�+��% `  ���@��t��%   =   tP�Å�t#�+��% `  ���@��t��%   =   t(�Å�t#�+��% `  ���@��t6��%   =   u(�E�P�E�Ph	�M��������7����M��E��M��E�o	���Ш�  �}� ��t#�+��% `  ���@��t4�}� ��t$�3�<@���	#�+����@��t�E�P�E�Ph�	�   �}� ��t#�+��% `  ���@��t4�}� ��t$�3�<����#�-   ���@��t�E�P�E�Ph�	�G�}� ��t#�+��% `  ���@��tF�}� tj ���X���	��#����@��t(�E�P�E�Ph�	�M��������#����M��E��M��E�}� ��t#�+��% `  ���@����t%   �%   ��t4�o	   u(�E�P�E�Ph�	�M��F�����������M��E��M��E���   t%�E�P�E�Ph�	�M������������E��M��E�E��M�H_^[�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���$SV�    W�5o	t0�%o	�����E�j P�_���	5o	YY�M܋E��M��H�!  �o	���?�   @�o	8u#8Hu�E�P�j����o	Y�@�o	�8 u�밍E�P�,����u�]�3�@Y��t��   t�E���e� ����#�:�~�E�0�X�  �o	� ����   <@��   �E�P�����E�Y����   �=o	 ��   �E�P�M��o	 �u�]�������o	�8@�u�]�u�]���   �E�P�I�����M�H�M���@�M�M�E��$d	�}����E�E܋E�E��E�P�M��m����u܋]��4�E܋E�hd	�M܉E��G����E܉E�E��E�E�P�M��7����u�]�]��u�}� t��t	��   �]�� �  ��tډ]���������   ��������o	� ��t<@t�E�`� ���  �@�X�o	�o	t)�}� u#��u�e� �e�  ���E�P�E�P����YY�p����E�P�u����YY���u��Mj�I����E_^[������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   SV�u3�W�� ���^!~��]�&  �o	� :��   <@�  8o	t8o	�]  9tSV�E�Phd	��p����S�����������E���E�F8]t'V�E�Pj[��h���������������E؉�E܉F�]�o	�9?�p  A�o	���$�I  H��   ��t^HH��   ��Vt��X���P��H���P� ���Y�>  �E�Pj]�E�PS�E�AjP�o	��������������������E�  �A�8_uK�y?uE�o	V��P���PS�E�SP�D���������������@�F�o	�8@��   �o	��   ��`���P�<���YP�E�Pj`�M�������������E�E��E�j'�M��E�����V�E�P�M��sj@ho	�M�����V�E�Ph	�M���������M����E���E�F��n	�9	tD�E�P�{����9��x���VIP�o	�E���E�VP�E�SjP����������������@�F8^������o	� :�t<@tJ!~�F��?9uj��������0V�E�Phd	�E�Pj�M��������������������@�F_��^[������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��o	���8��u�uj�u�����E���À�6|��9~��_t�E�`� ���  �@��S�ك�6@�o	��)u4���t�ك�=@�o	��|&����uj�u�I����E���L  ��x��~������u�E�`� ���  �@�%  �e� �e�  ��V�u�W�E��F�����E���   �E�P�E�Phd	�M��i�����������E�E��E�E��o	�8 tC�E�P�����YP�E�Pj �M�������������E��E�E�E�E�P�M��0����E�E��E��"�E�P�E�Pj�M���������r����E��E��E�E��o	� ����   <@��   �o	�o	��`<`�E�Ptq�[���Y��@�M��E�����   �o	���Ш�E�P��   ����YP�E�Pj �M��4�����������E��E�E�E�E�P�M��p����E�E��E�E��S�����YP�M������돋E�`� ���  �@�  �E�P�u�M�j������������~  ����YP�M������o	���Шt&�E�P�E�P�E�P�����Y���O�����@�M��E���E�P����YP�M��O���3�9t;�E�P�E�Pj(�M��V����������E��E�E�j)�M�E��:����E�E��E�E�Sj��n	�E���;�t�X�`� ������3��E�VP�s����E�P������P�E�Pj(�M�������������E��E�E�j)�M�E�������E�P�M������o	��`<`t;�t�E�P�M�������o	���Ш�E�Pt�����YP�M������������YP�M��O���;�t�E���E��F�M؋E��M܉H��Mj�k����E_^[��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���T�o	� SV�  ��!u�W3��E� ����  <$u.�u�E�P�EP�E�P�Y����Mԃ�;�t�E��M؉H�@  �o	�3�<A��!u��؉}�J��+��+�3�!u�U�Ã���   HtN���n  �o	���Ш��   ��t)�E�j �MԉUԉE�����j	������P�E��M��   j	�   �o	���Ш��   ��t7�E�j �M܉}܉E��@���j
�>�����P�E�P�M��R����8�@�}�E��j
������P�M������}��g�o	��������tW���ШtN��t7�E�j �M�U�E������j�������P�E��M�P�������@�M�E��j������P�M��@����o	�o	�8$u�u�E�P�EP�E�P������M̃���u#�o	�3�<A����J��+��+ڋU������E��M��J����9 tA�o	����   �uV�M��\���3��E܋EȉE��E�P�M��a����}� �E܋M��E�M�t4�M�j �M܉E�������E܉EԋE��E؍E�P�M��'����EԉE�E؉E���t7�E�j �Mԉ}ԉE������EԉE܋E؉E��E�P�M�������E܉E�E��E�����   �} t�E�`� ���  �@�  �> tx�E�P�E�Phd	�M�������� ����EĉE�EȉE��o	�8 �E�Pt�E�P�E�P����Y���������@�M���E�Pj�M������������EĉE�EȉE���o	�8 t�E�P�����YP�M������o	� ��uj�M�������o	<@�+����o	���Ш��t7��<uJ�} �����E�P�E�P�E�P�����Y���)�����@�M�E����<u�E�P����YP�M��"�����t(�E�P�E�Ph 	�M��f�����������EĉE�EȉE���t(�E�P�E�Ph�	�M��9����������EĉE�EȉE�3һ   9U��   �u9t`�N��uB�E9t;P�E�Pj �M��������m����EĉEԋE�j �MԉE�����V�E�P�M��J����7��   t��E���E��,V��E9t"P�E�Pj �M��Z����������E�P�M������M�ˀ}� t��    �E�U��5���9}uk�u9>tZ�F   uA�E98t:P�E�Pj�M��$����������EĉEԋE�j �MԉE������V�u�M������$Vj�u�z�������E98tP��Mj������E_^[������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� �E��  ��!U�3�!M�#o	��tq�:?u]�B<@u2�o	�E�P�Q���YP�E�Ph	�M��,����������M��E��3<$u �E�j P����YY��@<u�o	�o	�E�P����Y��@<u3���<t�o	   u�o	�: u�M��E���5o	�M������o	��u(�M���t��@�o	�����P��n	Y�o	��t>�5o	�M�P�����o	����� u@�
B�@�8 t���
B@���u����o	��������������������������������������������������������������������������������̋�U��QQ�o	� S3�V:���   <6|<9~<_uN�u�M�������E�u9t9t	�F   u	P�M�����9t	V�M������E�P�u����YY�E�   �uS�u�E�V�uP�v���3��>*��P�E�P�u趽���� ��j�M��,����u�M��N����u9t	V�M��F���W�}9t9t
j �M������W�M��'����M��E��M��H_^[���������������������������������������������������������������̋�U��h��u�u�u������E��]��������̋�U��hR��u�u�u�����E��]��������̋�U���u�u�u�u�����E��]��������jdhx*	�����}3�;�u3��rj�Ļ��Y��t�j�Q���Y�u��=�n	�E��n	�5�n	�5�n	�5�n	�EPV�u�u�u�M�������M�������E��n	�����E������	   �E�������j����Y���������������������������������������jdh�*	������}3�;�u3��rj����Y��t�j����Y�u��=�n	�E��n	�5�n	�5�n	�5�n	�u �u�u�u�u�M������M������E��n	�B����E������	   �E��8����j�����Y��������������������������������������̋�U��o	� ��$SVW���l  �o	�e� ���  ��!u��ǃ���E� ��NR�-  ��C��
�  ��-�$�h�	��  h�	��  h�	��  h�	��  h�	�  ��O��  ��  ��S��  ��X��  ��_��  �o	� �o	�E�����M��   ��L��   ��Ge��F}V��t=��$t�������   h�	�C  �u�E�P�g���Ph�	�u�������m  �o	j�M��.����H  h�	�  ��H|x��I~��Knh�	��   h�	��   ht	��   ��N��   ��OtW��RtK��Wt?�����w0�E��o	P�s����PY��M�U�����   �E��P��  hh	�~h\	�whP	�pj�[�E��e� !u��M�H�M�����4  hR��E�P�E�P�E�   	u�P��������u�uh$��M������M�E��M���   hH	�h� 	�M�������2�߃��"�E��5���hd 	�M�����h@	�M��\�������W����ǃ�Ct@jY+�t*+�t&+�t"+�t��uP�E���Et+�t+�t+�t+�u7�E�P�E�PhX 	��E�P�E�Ph4	�M��������^����E�E�E�E��E�8 t"P�E�Pj �M��z������4����E�P�M��¼���M�E��M��H�j�8 u8��t!h,	�M��������t!h 	�M��������th	�M�����h��E�P�E�P�u��������uj�u�������E_^[�Ë��	�	�	�	�	�   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����o	� S3۹  ��!M�+�V�]��s  ��$tj���ut.HtV�u����YY�c  h	�M��#���9t
j �M��r���h����v�o	�E��E�P�E�P�u��   �u���������  �o	�@<$t:���   �E�`� ���@���   �o	�o	� �u��Qp��   +�tc��AtJHt4Hu��o	!M�S�E�PhR��E�VP�]�����P�u�������   �o	jV�u�G����x�o	V�u�Z��������V�W��Rt*HtH�U����M�o	h�	課���@�o	�5���h	�M������9t
j �M��D���h��������uj�u��������E^[�������������������������������������������������������������������������������������������������������������̋�U����u�M�������o	� 3�:���   <?tG<Xt�E�P�u�;���YY�   �o	9M�u�Mh� 	螱���q�E�P�u�M�h	舱���T�o	�e�  ��Q�E�PhR��E�P�E�P�M��l�����M��@�E��E�P�u�Ƶ������E�P�u�M�j������譶���E����������������������������������������������������̋�U���Vj j��n	�������t�  �@ �`� �����3�V�u�����E�P�ڰ���E����E��E�j �M��E��[����u�E�P�M��������@�F�E^����������������������������������SVW�T$�D$�L$URPQQhpd�5    �B	3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C������   �C�����d�    ��_^[ËL$�A   �   t3�D$�H3��>���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�!���3�3�3�3�3���U��SVWj RhQ����_^[]�U�l$RQ�t$������]� ����������������������������������������������������������������������������������������������U��W�}3�������ك��E���8t3�����_������������̋�U����u�M������E����   ~�E�Ph  �u�O���������   �M�H%  �}� t�M��ap�����������������������̋�U��=�o	 u�E��N	�A%  ]�j �u����YY]������������̋�U����u�M��n����E����   ~�E�Pj�u����������   �M�H���}� t�M��ap����������������������̋�U��=�o	 u�E��N	�A��]�j �u誷��YY]�����������̋�U����u�M�������E����   ~�E�Pj�u����������   �M�H���}� t�M��ap����������������������̋�U��=�o	 u�E��N	�A��]�j �u�����YY]�����������̋�U����u�M��2����E����   ~�E�Pj�u�o���������   �M�H���}� t�M��ap����������������������̋�U��=�o	 u�E��N	�A��]�j �u�$���YY]�����������̋�U����u�M������E����   ~�E�Ph�   �u�����������   �M�H%�   �}� t�M��ap�����������������������̋�U��=�o	 u�E��N	�A%�   ]�j �u荾��YY]������������̋�U����u�M�������E����   ~�E�Pj�u�*���������   �M�H���}� t�M��ap����������������������̋�U��=�o	 u�E��N	�A��]�j �u�{���YY]�����������̋�U����u�M��O����E����   ~�E�Pj�u����������   �M�H���}� t�M��ap����������������������̋�U��=�o	 u�E��N	�A��]�j �u�|���YY]�����������̋�U����u�M������E����   ~�E�Ph  �u�����������   �M�H%  �}� t�M��ap�����������������������̋�U��=�o	 u�E��N	�A%  ]�j �u����YY]������������̋�U����u�M��
����E����   ~�E�PhW  �u�D���������   �M�H%W  �}� t�M��ap�����������������������̋�U��=�o	 u�E��N	�A%W  ]�j �u�%���YY]������������̋�U����u�M��c����E����   ~�E�Ph  �u����������   �M�H%  �}� t�M��ap�����������������������̋�U��=�o	 u�E��N	�A%  ]�j �u�~���YY]������������̋�U����u�M�輿���E����   ~�E�Pj �u�����������   �M�H�� �}� t�M��ap����������������������̋�U��=�o	 u�E��N	�A�� ]�j �u����YY]�����������̋�U��}�   ���]����̋�U��E��]���̋�U���u�u����YY��u�}_t]�3�@]��������̋�U���u�,���Y��u�}_t]�3�@]�������̋�U���u�u����YY��u�}_t]�3�@]��������̋�U���EP�
���Y��u�}_t]�3�@]��������̋�U��E�� ]���̋�U���SV�u�M��A����]�   ;�sT�M胹�   ~�E�PjS�t����M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P蓯��YY��t�Ej�E��]��E� Y������ *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�=�����$���o������E�t	�M�����}� t�M��ap�^[����������������������������������������������������������������������̋�U��=�o	 u�E�H���w�� ]�j �u�����YY]�����������̋�U���(�B	3ŉE�SV�uW�u�}�M�蟼���E�P3�SSSSW�E�P�E�P�O����E�E�VP������(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������������������������������������������������̋�U��j �u�u�=�����]�����̋�U���(�B	3ŉE�SV�uW�u�}�M�豻���E�P3�SSSjW�E�P�E�P�`����E�E�VP������(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�����������������������������������������������̋�U��j �u�u蹷����]�����̋�U���(�B	3ŉE�SV�uW�u�}�M��º���E�P3�SSSSW�E�P�E�P�r����E�E�VP�P�����(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[� ����������������������������������������������̋�U��j �u�u������]�����̋�U��EV�5lo	�����t������    �y�����lo	��^]������������̡lo	Ë�U��MS�YV�u3�;�u����j^�0�6������   9Ev�U�;�~��@9Ew�e���j"Y�����W�~�0�ǅ�~���t��C�j0Y�@J���M�  ��x�;5|�� 0H�89t�� �>1u�A�W蚭��@PWV�_�����3�_^[]��������������������������������������������̋�U��Q�M�AS����% �  V��  #�W�E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��B��<  �U����������U��E����������Ɂ���  ��P��t�M�_^f�H[���������������������������������������������̋�U���0�B	3ŉE��ES�]V�E�W�EP�E�P�%���YY�E�Pj j���uЋ���f��D����u܉C�E��E��C�E�P�uV�������$��u�M�_�s^��3�[�W�����3�PPPPP�)����������������������������������������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ����������������������������������������������������������������̀�@s�� s����Ë�3Ҁ����3�3���������j�����Y��̋�U��E�M%����#�V�u������t$��tj j 腤��YY�����j^�0�V������P�u��t	�a������X���YY3�^]�����������������������̋�U��M��tj�3�X��;Es�R����    3�]��MV���uF3����wVj�5a	���	��u2�=xh	 tV�n���Y��uҋE��t�    3���M��t�   ^]��������������������������������̋�U��} u�u�R���Y]�V�u��u�u�l���Y3��MW�0��uFV�uj �5a	���	����u^9xh	t@V�ϸ��Y��t���v�V迸��Y�^����    3�_^]��M�������	P�V���Y����5�������	P�>���Y�����������������������������������������������̋�U��MS3�;�vj�3�X��;Es������    3��A�MVW��9]t�u脳��Y��V�u������YY��t;�s+�Vj �S��������_^[]����������������������������jh�*	�0����°���@x��t�e� ���3�@Ëe��E�����������˷�����������������臰���@|��t��鈦������jh�*	�Һ���5po	�ԑ	��t�e� ���3�@Ëe��E������M������������������h\��ܑ	�po	����̋�U��E�to	�xo	�|o	��o	]��������jh�*	�R���3�W����Y�}�9}u�to	�5to	�ԑ	�E��E�   ��xo	�5xo	�ԑ	�E��E�   ;�t��t�7�����E������   9}�u3��3�W�p���YÃ}�t�u��U�Y3�@茶��� ��������������������������������������̋�U��E�\�V9Pt��k�u��;�r�k�M^;�s9Pt3�]���������������5|o	�ԑ	�����ٮ����d����ή����`���jh+	�%����e� �u�]����  ����  j_;���   ����   ����   ����   ����   ��t��t	����  �c���������  ���9~\u'�5X�膙��Y�F\���t  �5X�WP�)������v\�������Y���Q  �H�M�M���.  ����H���\�k�V\�x�;��  9t��  j ����Y�e� ;�t��u>�=�o	 u5jhX'���	3�A;�u��o	����������	��E�   �u��+�ty��t��	tN��t(H��   �5|o	�ԑ	�E�;�toV�ܑ	�|o	�a�5xo	�ԑ	�E�;�tNV�ܑ	�xo	�@�5�o	�ԑ	�E�;�t-V�ܑ	��o	��5to	�ԑ	�E�;�tV�ܑ	�to	�E������   �}� u�E��8�]j 蹴��YÃ�t$��t��t��~��~�5����    ��������蹳���������������������������������������������������������������������������������������������������������������������������������������������������j h8+	�U���3��}�}؋]��Kt��jY+�t"+�t+�tY+�uC�ʗ�����}؅�u����T  �to	�to	�U�w\���g���Y�p��Q�Ã�t2��t!Ht�����    ����빾|o	�|o	��xo	�xo	�
��o	��o	�E�   P�ԑ	�E�3��}���   9E�uj脡��9E�tP�?���Y3��E���t
��t��u�O`�MԉG`��u>�Od�M��Gd�   ��u,�P��M܋T�P�9M�}�M�k��W\�D�E����Y�����E������   ��u�wdS�U�Y��]�}؃}� tj 聲��Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3�膱����������������������������������������������������������������������������������������������������������̋�U��E��o	]���̋�U��QV�5�o	�ԑ	���E��u�S���j^�0��������   �  W����   h	���	�E���u����j^�0��������   h�	P� �	����u(������5�	����P�����Y�������P����Y�LSV�ܑ	���Ѥ��Wh�o	�����	;�[t	�u����	j�u�օ�u虿���    莿��� �3�_^���������������������������������������������������������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]���������������������������̋�U��E�H<��ASV�q3�W�D��t�}�H;�r	�X�;�r
B��(;�r�3�_^[]����������������������������̋�U��j�hX+	h��d�    P��SVW�B	1E�3�P�E�d�    �e��E�    h   �x�������tT�E-   Ph   �+�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE�3ҁ9  ���Ëe��E�����3��M�d�    Y_^[��]�����������������������������������������������̋�U����u�M�袩���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap����������������������̋�U��jj �u�u������]������̋�U��jj �uj �g�����]������̋�U��jj �u�u�H�����]������̋�U��jj �uj �*�����]������̋�U��jj �u�u������]������̋�U��jj �uj �������]������̋�U��jh  �u�u�������]�������̋�U��jh  �uj ������]������̋�U��jh  �u�u������]�������̋�U��jh  �uj �e�����]������̋�U��jh  �u�u�C�����]�������̋�U��jh  �uj �!�����]������̋�U��jhW  �u�u�������]�������̋�U��jhW  �uj �������]������̋�U��jj�u�u������]������̋�U��jj�uj ������]������̋�U��jj �u�u������]������̋�U��jj �uj �c�����]������̋�U��jj �u�u�D�����]������̋�U��jj �uj �&�����]������̋�U����u�M�车���E��t*�x�  u!jj �u�u��������}� t�M��ap��À}� t�E��`p�3�����������������������̋�U��j �u�A���YY]����̋�S��QQ�����U�k�l$���   �B	3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����$�������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P������h��  ��x���������>YYt�= Q	 uV����Y��u�6�����Y�M�_3�^�������]��[�������������������������������������������������������������������������������̋�U���$�B	3ŉE��ES�E��EVW�E�蝝���e� �=�o	 �E�u}h�	���	�؅��  �= �	h�	S�ׅ���   �5ܑ	P��hx	S��o	��P��h`	S��o	��P��h@	S��o	��P�֣�o	��th$	S��P�֣�o	��o	�M�5ԑ	;�tG9�o	t?P���5�o	���֋؅�t,��t(�ׅ�t�M�Qj�M�QjP�Ӆ�t�E�u	�M    �3��o	;E�t)P�օ�t"�ЉE��t��o	;E�tP�օ�t�u��ЉE��5�o	�օ�t�u�u��u��u����3��M�_^3�[�5�����������������������������������������������������������������������������������������������̋�U��V�uW��t�}��u�ֶ��j^�0�{�����_^]ËM��u3�f��݋�f�: t��Ou��t�+��f�
��f��tOu�3���u�f�脶��j"Y��������������������������������̋�U��US�]VW��u��u9Uu3�_^[]Å�t�}��u�,���j^�0�Ѷ�����݅�u3�f��ЋM��u3�f��ԋ��u��+��f���f��t'Ou��"��+��f���f��tOtKu��u3�f����y���3����u�MjPf�DJ�X�d���f�蝵��j"Y����j�����������������������������������������������������̋�U��Ef���f��u�+E��H]������̋�U��V�uW��t�}��u�#���j^�0�ȵ����_^]ËE��uf��ߋ�+��f���f��tOu�3���u�f�����j"Y���������������������������̋�U��M��x��~��u�\_	]á\_	�\_	]�蓴���    �7������]���������������̋�U��E�`_	]����3�Ë�U��QQ�E���]��E�������̃%$�	 ��̋�U��ES3�VW9]u;�u9]u3�_^[]�;�t�};�w�
���j^�0说������9]u��ҋU;�u��ك}���u��+�
�B:�t"Ou����+���A:�tOt�Mu�9]u�;�u��}�u�MjP�\�X�x����萳��j"Y������������������������������������������������̋�U����B	3ŉE��E� �@SVW�=��	3�VV�u�E��u�׋ȉM�;�u3��   ~Ej�3�X���r9�D	=   w�5�����;�t����  ���P�{���Y;�t	� ��  �����3�;�t��u�S�u�u�ׅ�t VV9uuVV��u�uj�SV�u��L�	��S�~���Y�ƍe�_^[�M�3��j����������������������������������������������������������̋�U����u�M��A����u�E��u�u�uP��������}� t�M��ap����������������̋�U��QQ�EV�u�E��EWV�E��������Y;�u�ױ��� 	   �ǋ��J�u�M�Q�u�P�Ē	�E�;�u��	��t	P�R���Y�ϋ�������	�����D0� ��E��U�_^�����������������������������������jhx+	� �������]܉]��E���u�����  �2���� 	   �Ë��   ��x;T�	r�����  �
���� 	   讱���ы����<���	��������L1��t�P�Q���Y�e� ��D0t�u�u�u�u萍�����E܉U��訰��� 	   �q����  �]܉]��E������   �E܋U�������u�����Y����������������������������������������������������������̋�U���  �����B	3ŉE��EV�uW3���4�����8�����0���9}u3��  ;�u����8�����    苰������  ������S����	������L8$�����$�����?�����t��u'�M����u�d����  舯���    �,����  �D8 tjj j V�=�����V�ק��Y����  ��D���  記���@l3�9H�� �����P��4���̒	3�;��`  ;�t8�?����P  �Ȓ	��4����� ���3���,���9E�#  ��@�����?������g  ���$���3���
��������ǃx8 t�P4�U�M��`8 j�E�P�K��P�#���Y��t:��4���+�M3�@;���  j��D���SP�ڈ���������  C��@����jS��D���P趈��������n  3�PPj�M�Qj��D���QP�� ���C��@����L�	�����=  j ��,���PV�E�P��$���� �4�l�	���
  ��@�����0������8���9�,�����  ����� ��   j ��,���Pj�E�P��$���� �E��4�l�	����  ��,�����  ��0�����8����   <t<u!�33Ƀ�
������@�����D��������<t<uR��D����Ŭ��Yf;�D����I  ��8�������� t)jXP��D���蘬��Yf;�D����  ��8�����0����E9�@���������  ����8����T4��D8��  3ɋ�D8���  ��?��� ��D�����   ��4���9M��  ��3�+�4�����H���;Ms&�CA�� �����
u��0���� @F�@F���  rՋ���H���+�j ��(���PV��H���P��$���� �4�l�	���C  ��(����8���;��;  ��+�4���;E�l����%  ��?�����   ��4���9M�H  ��@��� ��+�4���j��H���^;MsC��Ή� �����
u�0���j[f��� �����@����@���f�Ɓ�@����  r�����H���+�j ��(���PV��H���P��$���� �4�l�	���i  ��(����8���;��a  ��+�4���;E�G����K  ��4�����,���9M�u  ��,�����@��� +�4���j��H���^;Ms;��,�����,���΃�
uj[f���@����@���f�Ɓ�@����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �L�	��;���   j ��(���P��+�P��5����P��$���� �4�l�	��t�(���;�����	��D���;�\��,���+�4�����8���;E�����?Q��(���Q�u��4����48�l�	��t��(�����D��� ��8������	��D�����8��� ul��D��� t-j^9�D���u詩��� 	   �r����0�?��D����>���Y�1��$���� �D@t��4����8u3��$�i����    �2����  ������8���+�0���[�M�_3�^�%��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������jh�+	�@����]���u�7����  �[���� 	   ����   ��x;T�	r�����  �4���� 	   �ا���ҋ����<���	�������D0��t�S�{}��Y�e� ��D0t�u�uS�}�����E���ڦ��� 	   裌���  �M���E������   �E��K���Ë]S�.}��Y�����������������������������������������������������̋�U����o	h   �{��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]������������������̋�U��E���u����� 	   3�]Å�x;T�	r����� 	   菦���ދȃ�������	���D��@]���������������������̸(Q	á �	Vj^��u�   �;�}�ƣ �	jP躧��YY��o	��ujV�5 �	衧��YY��o	��ujX^�3ҹ(Q	���o	��� �����S	|�j�^3ҹ8Q	W��������	����������t;�t��u�1�� B���Q	|�_3�^���������������������������������������������褄���=�_	 t�ԇ���5�o	�q���Y��������̋�U��V�u�(Q	;�r"���S	w��+�����Q�����N �  Y�
�� V���	^]����������������̋�U��E��}��P�ǁ���E�H �  Y]ËE�� P���	]������������̋�U��E�(Q	;�r=�S	w�`���+�����P�J���Y]Ã� P���	]���������������̋�U��M�E��}�`�����Q����Y]Ã� P���	]�����������̋�U��E��u�}����    �!������]Ë@]����������jh�+	�#���3�3�9u��;�u�@����    ��������_�ܒ��j [�Pj�ڥ��YY�u��Œ���P��}��Y���EPV�u譒���P�����E�蝒���PW�<������E������	   �E��c�����w����� Pj�Ɨ��YY�����������������������������������������̋�U��EP�u�u�%v����]������̋�U��EP�u�u襆����]������̋�U��EPj �u臆����]������̋�U��EP�u�u�w�����]������̋�U��EPj �u�Y�����]������̋�U��B	�U��3�9�o	�����#щ�o	]����������̡B	��3�9�o	���������̋�U���SV�u3�W�};�u;�v�E;�t�3��{�E;�t�������v�h���j^�0�������V�u�M��Y����E�9X��   f�E��   f;�v6;�t;�vWSV�}��������� *   ����� 8]�t�M��ap�_^[��;�t&;�w ����j"^�0藡��8]�t��E��`p��y�����E;�t�    8]��<����E��`p��0����MQSWVj�MQS�]�p�L�	;�t9]�j����M;�t�����	��z�P���;��s���;��k���WSV��|�����[���������������������������������������������������������������������������������������̋�U��j �u�u�u�u虇����]�������̋�U����u�M���M��̋���E�P�u�E����   �E��uP�Z�������u�E������}� t�M�ap����������������������̋�U��Q�M��j �u诛��P�u�E�P��������u�E��Ã����������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ������������������������������������̋�U��M�I�8 t@��u�I�E+�H]�������̋�U����B	3ŉE��US3�VW;�~�E��I8t@;�u������+�H;�}@�E�]�9]$u�E� �@�E$�5Ԓ	3�9](SS�u���u��   P�u$�֋��}�;�u3��R  ~Cj�3�X����r7�D?=   w������;�t� ��  �P�:~��Y;�t	� ��  ���E���]�9]�t�W�u��u�uj�u$�օ���   �5В	SSW�u��u�u�։E�;���   �   �Mt)�E ;���   9E���   P�uW�u��u�u���   �}�;�~Bj�3�X����r6�D?;�w�7�����;�th���  ���P�}}��Y;�t	� ��  �����3�;�t?�u�W�u��u��u�u�օ�t"SS9] uSS��u �u�u�WS�u$�L�	�E�W�x���Y�u��o����E�Y�e�_^[�M�3��Z�����������������������������������������������������������������������������������������������������������������������������̋�U����u�M������u(�E��u$�u �u�u�u�u�uP�l�����$�}� t�M��ap�������������������̋�U��QQ�B	3ŉE�S3�VW�]�9]u�E� �@�E�5Ԓ	3�9] SS�u���u��   P�u�֋�;�u3��~<�����w4�D?=   w�k~����;�t� ��  �P�{��Y;�t	� ��  ���؅�t��?Pj S�w����WS�u�uj�u�օ�t�uPS�u�ؒ	�E�S踘���E�Y�e�_^[�M�3�裞������������������������������������������������������������̋�U����u�M��w����u$�E��u�u�u�u�uP�������}� t�M��ap������������������̋�U���S�XBV���HD�M���u�����  �e� W�E�FPj1S�E�jP��{�����FPj2S�E�jP��{����FPj3S�E�jP�{����FPj4S�E�jP�{����P��FPj5S�E�jP�{����FPj6S�E�jP�x{��Vj7S��E�jP�g{����F Pj*S�E�jP�S{����P��F$Pj+Sj�E�P�<{����F(Pj,S�E�jP�({����F,Pj-S�E�jP�{����F0Pj.S�E�jP� {����P��F4Pj/S�E�jP��z����FPj0S�E�jP��z����F8PjDS�E�jP��z����F<PjES�E�jP�z����P��F@PjFS�E�jP�z����FDPjGS�E�jP�z����FHPjHS�E�jP�nz����FLPjIS�E�jP�Zz����P��FPPjJS�E�jP�Cz����FTPjKS�E�jP�/z����FXPjLS�E�jP�z����F\PjMS�E�jP�z����P��F`PjNS�E�jP��y����FdPjOS�E�jP��y����FhPj8S�E�jP��y����FlPj9S�E�jP�y����P��FpPj:S�E�jP�y����FtPj;S�E�jP�y����FxPj<S�E�jP�uy����F|Pj=S�E�jP�ay����P����   Pj>S�E�jP�Gy������   Pj?S�E�jP�0y������   Pj@S�E�jP�y������   PjAS�E�jP�y����P����   PjBS�E�jP��x������   PjCS�E�jP��x������   Pj(S�E�jP�x������   Pj)S�E�jP�x����P����   Pj�u��E�jP�x������   Pj �u��E�jP�nx������   Ph  �u��E�jP�Rx������   Ph	  �u��E�j P�6x����E���P���   ���   Pj1S�E�jP�x������   Pj2S�E�jP��w������   Pj3S�E�jP��w������   Pj4S�E�jP��w����P����   Pj5S�E�jP�w������   Pj6S�E�jP�w������   Pj7S�E�jP�w������   Pj*S�E�jP�ow����P����   Pj+S�E�jP�Uw������   Pj,S�E�jP�>w������   Pj-S�E�jP�'w������   Pj.S�E�jP�w����P����   Pj/S�E�jP��v������   Pj0S�E�jP��v������   PjDS�E�jP��v������   PjES�E�jP�v����P����   PjFS�E�jP�v������   PjGS�E�jP�v�����   PjHS�E�jP�iv�����  PjIS�E�jP�Rv����P���  PjJS�E�jP�8v�����  PjKS�E�jP�!v�����  PjLS�E�jP�
v�����  PjMS�E�jP��u����P���  PjNS�E�jP��u�����  PjOSj�E�P��u�����   Pj8S�E�jP�u�����$  Pj9S�E�jP�u����P���(  Pj:S�E�jP�zu�����,  Pj;S�E�jP�cu�����0  Pj<S�E�jP�Lu�����4  Pj=S�E�jP�5u����P���8  Pj>S�E�jP�u�����<  Pj?S�E�jP�u�����@  Pj@S�E�jP��t�����D  PjAS�E�jP��t����P���H  PjBS�E�jP�t�����L  PjCS�E�jP�t�����P  Pj(S�E�jP�t�����T  Pj)Sj[�E�SP�ut����P���X  Pj�u��E�SP�Zt�����\  Pj �u��E�SP�Bt����`  Vh  �u���E�SP�'t����<�_^[��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��V�u���c  �v�ގ���v�֎���v�Ύ���v�Ǝ���v辎���v趎���6诎���v 觎���v$蟎���v(藎���v,菎���v0臎���v4�����v�w����v8�o����v<�g�����@�v@�\����vD�T����vH�L����vL�D����vP�<����vT�4����vX�,����v\�$����v`�����vd�����vh�����vl�����vp������vt�����vx�����v|������@���   �֍�����   �ˍ�����   ��������   赍�����   認�����   蟍�����   蔍�����   艍�����   �~������   �s������   �h������   �]������   �R������   �G������   �<������   �1�����@���   �#������   �������   �������   �������   ��������   �������   �������   �֌�����   �ˌ�����   ��������   赌�����   誌�����   蟌����   蔌����  艌����  �~�����@��  �p�����  �e�����  �Z�����  �O�����  �D�����   �9�����$  �.�����(  �#�����,  ������0  ������4  ������8  �������<  ������@  ������D  �֋����H  �ˋ����@��L  轋����P  貋����T  觋����X  蜋����\  葋����`  膋����^]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��SV�u�~  W� L	tBhd  j�������YY��u3�@�I�Ƌ��v�����tW����W�[���YY��Ǉ�      ������   ;�t�   P��	���   3�_^[]��������������������������������2�8tSV�<0|<9,0�A8u�^[�<;u���X�@8u��������������̋�U��V�u��tY�;8T	tP讉��Y�F;<T	tP蜉��Y�F;@T	tP芉��Y�F0;hT	tP�x���Y�v4;5lT	tV�f���Y^]��������������������������̋�U���SV�uW3��u��}�9~u9~u�}��}��8T	�e  jPj脌����YY;�u3�@�  ���   jY��j���^��3�Y�E�;�u	S�ۈ��Y�ыu�89~��   j�^��Y�E�;�u3�FS貈���u�誈��YY���D  �8�v>SjV�E�jP�k�����CPjV�E�jP�k����CPjV�E�jP�k����C0PjV�E�jP�wk����P��C4PjV�E�jP�`k�����tS����Y����k����C����0|��9��0�@�8 u��>��;u���N�F�> u���8T	��<T	�C�@T	�C�hT	�C0�lT	�}��C4�M��u3�@��M���t����   �=�	��tP�׋��   ��tP�ׅ�u���   脇�����   �y���YY�E����   �E����   ���   3�_^[������������������������������������������������������������������������������������������������������������������������������2�8tSV�<0|<9,0�A8u�^[�<;u���X�@8u��������������̋�U��V�u����   �F;DT	tP�~���Y�F;HT	tP�l���Y�F;LT	tP�Z���Y�F;PT	tP�H���Y�F;TT	tP�6���Y�F ;XT	tP�$���Y�F$;\T	tP����Y�F8;pT	tP� ���Y�F<;tT	tP����Y�F@;xT	tP�܅��Y�FD;|T	tP�ʅ��Y�FH;�T	tP踅��Y�vL;5�T	tV覅��Y^]���������������������������������������������������������������̋�U���SV�uW3��}��u��}�9~u9~u�}��}��8T	��  jPj蜈����YY;�u3�@�  j��Z��Y�E�;�u	S����Y���89~�4  j��Z��Y�E�;�uS�߄���u��ׄ��Y�҉8�v8�CPjV�E�jP��g�����CPjV�E�jP��g����CPjV�E�jP�g����CPjV�E�jP�g����P��CPjV�E�jP�g����C PjPV�E�jP�|g����C$PjQV�E�jP�hg����C(PjV�E�j P�Tg����P��C)PjVj �E�P�=g����C*PjTV�E�j P�)g����C+PjUV�E�j P�g����C,PjVV�E�j P�g����P��C-PjWV�E�j P��f����C.PjRV�E�j P��f����C/PjSV�E�j P��f����C8PjV�E�jP�f����P��C<PjV�E�jP�f����C@PjV�E�jP�f����CDPjV�E�jP�of����CHPjPV�E�jP�[f����P��CLPjQV�E�jP�Df�����t$S�}��S�
����u������u��������������C����0|��9��0�@�8 u�� ��;u���N�F�> u���jY�8T	���E���   �	����   �I�u�K���   �I�K���   �I0�K0���   �@4�M��C43�@3��9}�t�M�����   ;�tP��	���   ;�t#P��	��u���   �/������   �$���YY�E����   �E����   ���   3�_^[����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������k���Hl;�N	t�L	�Hpu�u����T	���������̡�T	��k���ȋAl;�N	t�L	�Qpu�]u�����   ����������̋�U��j
j �u��b����]�����̋�U���uj
j �u�e����]������̋�U��]�����̋�U��]��f���̋�U��j
j �u�[����]�����̋�U���uj
j �u�x����]������̋�U��=��	 V�5�_	u3��cW��u95�_	tS��T����uJ�5�_	��t@�} t:�u�a��Y���'P�a��Y;�v��<8=uW�uP�it������t�����u�3�_^]Ë�D8����������������������������������̋�U��SV��3�;�u贀��j^�0�Y������C�E�;�t9]w��9]u�;�t�W�u�GW����Y;�t/W�a��@Y�9]t ;Evj"X_^[]�W�u�u�Ł������u3���SSSSS�w������������������������������������̋�U��VW��3�;�u����j^�0謀�����O�E�7;�t�09ut�S�u�V����Y;�tKS�a`���pjV�[`���3���;�u����    ���� [_^]�SVP��������u�E;�t�03���WWWWW�Hv������������������������������������������jh�+	�s��3�9E����u�;���    ����3��?��  V�u��t��YY;����t�j�\��Y�e� �u��U��Y�E��E������	   �E��o���j�Dp��Y�������������������������������jh�+	�r��j�9\��Y3ۉ]�3��};���;�u�~��j^�0�9���u��j��M;�t	9]w	;�u
9]u3�@�3�;�t�;�t��u�U��Y��;�t0V��^��Y@�9]t!;Ev	�E�"   �V�u�u�����;�u�]��E������   �E��n���SSSSS��t��j�Yo��Y����������������������������������������������������jh,	�q��j�9[��Y3��u�3��};���;�u�}��j^�0�9~���u��t�7�E;�t�03�9u��;�t��u�+T��Y��;�t�S��]���pjV��]�����3�;�u�>}���    �3}��� �E��SVP�~����;�u!�E;�t�0�}��E������   �E��m���WWWWW�s��j�On��Y�����������������������������������������������������̋�U���L�B	3ŉE�S3�V�uW�]ԉ]�]��]؉]܉u��]�9^�  �F9u P�F0h  P�E�SP�L^��������  j�Q��j��  W�E��x~��jW�E��m~��jW�E��b~��jh  �E��S~����$�E�9]��  9]��v  ;��n  9]��e  9]��\  �Eԉ3��M܈@=   |�E�P�v���	���2  �}��(  �E�EЃ�~.8]�t)�E�:�t �x�����M�� �G;�~��8X�uڋE�SS�v   Ph   �u܉E�jS��j���� ����  �M��E�S�v��   W���   QW@Ph   �vS��k����$����  �E�S�v�   WP�E�W@Ph   �vS��k����$���b  �E�}����   3҃}�f��U؉Mč��   �_�Z��M����   �MȈ~U8]�tP�M�M�:�tD�I��҉M�;�(��H   ��M��E� �  f����M̋M��	9M�~�M���M�8Y�u�h�   ��   QP�e��j��   PW�e���E�j��   QP�e�����   ��$;�tKP��	��u@���   -�   P��x�����   ��   +�P�x�����   +�P�x�����   �x�����E��    ���   �E����   �Eĉ��   �E����   �Eȉ��   �EЉ��   �u��Ux��Y���o�u��Hx���u��@x���u��8x���u��0x��3ۃ�C�ˋ��   ;�tP��	���   ���   ǆ�   �	ǆ�   @
	ǆ�   �	ǆ�      3��M�_^3�[��|����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������a���ȋAl;�N	t�L	�Qpu�Pk�����   ����������̋�U��E��u]�.t��� ���   ]���������0a���ȋAl;�N	t�L	�Qpu��j���@�����������a���ȋAl;�N	t�L	�Qpu��j���@������������`���ȋAl;�N	t�L	�Qpu�j�������������̡�o	ø�o	Ë�V���t��t;�tWj6Y���  P�~p��Y_^���������̋�U��V�b`���Hpj Z���r�U���t0��t3��t��t��v���    �uw�������������Hp��L	���^]�����������������������̡�N	���   ��T	���   ��T	���   ��U	�����������jh8,	�"j���u����   j��S��Y�e� �F��tP��	��u�F=�E	tP��t��Y�E������[   �> t<j�S��Y�E�   �6�`p��Y���t�8 u=�M	tP�({��Y�E������&   �𭺉�FV�t��Y�Lf��Ëuj�g��YËuj�g��Y������������������������������������������������̋�U��]��S����jhh,	�#i���^����jj�}w��YY���u��u�3u���    3��[�rh����k���Gl��Gh�Fj�R��Y�e� �6�ln��Y�E������/   j�yR��Y�E�   �v��	�E������   ���`e��Ëu�j�"f��YËu�j�f��Y���������������������������������������������zk��3�Ë�U��SW3�3�9]~"V�u���6�u�u�F������uG;}|�^_[]�SSSSS�k������������������̋�U��SVW�}h�   3�SW�P���u�����u3���   <.u1�F8t*jP���   jP��K������u���   ��SSSSS�j��h�	V�]��E��;��   �} �<0�u��@��   ��.t|PVj@�u�;�}u��@sh��_tcP�EVj@��@��}uQ��sL��t��,uCP�EVj��P�^K������u4��,�=������5����E�wh�	V�OE����YY�k������_^[]�3�PPPPP�=�������������������������������������������������������������������������̋�U��SV�uV�u�u�"t����3ۅ�uA�F@8tPh�	j�u�u�~E�������   8^[tPh�	j�u�u�\E����]�SSSSS�$i����������������������������̋�U���S3�ChU  �]���F��Y�E����=  W�x� ��vX�Q  h<��5�	jSW��D���FX���E��	�E�h�	SW�1D��������   �E��H�1�M��0�R��YY��t�e� �E��0�E�h<��E��E��0jSW�D�����}��	|��}� uU�FP��	��tP�Ӆ�u	�vP�,p��Y�FT��tP�Ӆ�u	�vT�p��Y�E��fT �fL �FP�~H���Z3�PPPPP��g���u���o���FP�=�	3�Y;�tP�ׅ�u	�vP��o��Y�FT;�tP�ׅ�u	�vT�o��Y�Fh�^T�^L�^P�^H_[������������������������������������������������������������������������������������������̋�U���   �B	3ŉE��ESV�uW�}��d����E��\�����`����Y�����   ��T������   ���   K  ��X�����h�������  ��d��� ��  �} ��  �>CuS�~ uMh�	�u��d����Tq������u'��tf�f�Gf�G��`�����t�  ��d����C  3�PPPPP�pf��V�0P����   Y��P���;�s,V��h����xP��YY����   V��X����bP��YY����   ��L��� ��l���VP�oM��YY����   ��l���PSP�O��������   �C��T������l���PW��h����oQ�����> t
��P���;�r��L����R�@PVW��X�����F�������%���3�9�\���tjS��\����0Z����9�`���tj��T�����`����Z������h����u��d�����o������u��h����VVVVV�����3��M�_^3�[�Lr�������������������������������������������������������������������������������������������������������������������������������������������̋�U����  �B	3ŉE��ES��W��p�����h����W����S��\���P��P���Ph�   ��x���P��h����h������u3��M�_3�[�Xq��������sH��x���P�LN��YY��u�CH�Ӎ�x���P��M����P��t�����A��YY��l�����t��CH��p�����h����D���X���� ��H����Ak��jP��d�����8���P�YX���F��x���Q��t�����L�����l��������QP�3n�������	  ��l�����X������CH��P����j��P���P��d�����W������p����  ��\�����t��� �F���  ���  ��d������  �V;t6���t������d�����@����P�H��@�������t�����d���|��-��t�����t#����  ����  �P���  ���d����H��t���urj�v��x����vPjh	jj �K[���� ��t<3���  f!�Ex���@��r�h�   �5(U	��x���P��V�������@���  ����   �F���  ���  ���   ��p���u	��\����F��p���k�V���	Y��t1��h�����l����CH��i����H���Y��X������L����F������h���L	t.��p�������4���	��u�4��i���sT�i���cL YY��p�����l�������    ���Y���3�PPPPP�ia����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���   �B	3ŉE��ESV3ۋ�W��h���;�t;�tP�����Y��  ɋD�H��  ǅp���   ��t���;���  �8L�0  �xC�&  �x_�  ��h�	W�<����YY����   +ǉ�p�����   �;;��   ǅl���   ��	���p���PW�6�^������u�6�I��Y9�p���t��l��������	~�Ch�	S��:����3�YY;�u	�;;��   ��l���DWS��x���h�   P�@������uT��l�����h�����=x�����x���P����Y��t��t�����? t
G�? ����3�9�t�����   ��h����   VVVVV�	_��3��xSSSh�   ��x���QP�Ac����;�t\�~H��t5�7��x���P��H��YY��t��x���P������Y��u!�p������t���C����~�3�9�p���u9�t���t�����M�_^3�[�k������������������������������������������������������������������������������������������������������������������������������������������̋�U��}VWw$�} t3�GWj�Ki����YY��u�g���    3�_^]�Wh�   �'i��YY���u	V�e��Y��Wh   �i��YY�F��u�6�e��V�e��Y�ً��M	�w����u�M������Y��u�6�a���6��k��V�Ke�����2�v��p��D��YY��t#�v�+e���6��`���6�k��V�e����3��
�F�8�F�8���>���������������������������������������������������������������̋�U��]��S����jh�,	�Y���e� �}v��e���    �yf��3��9  �%O�����u��Y���Np�e� 3�GWh�   ��g��YY�؉]܅���   j�C��Y�}��Nl���E����e� �   �u�M������Y�E�����   �} thL	�u�7F��YY��t�=�o	j�B��Y�E�   �~lSW�$a��S�_�����Fpu?�L	u6�7h�N	� a��YY��N	���   ��T	���   ��T	���   ��U	�e� �   �.�]܋u�3�Gj�V��YËu�j�V��Y��S�_��S��i��YY�E������   �E��U��Ëu�fp����������������������������������������������������������������������������������������������̋�U��Q���  f9Eu3��ø   f9Es�E��T	�A��E�Pj�EPj�ؒ	��u!E��E��M#�����������������������̋�U��]�P���̋�U���u�u�P��YY]���������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ����������������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ����������������������������U��SVWUj j h��u�P��]_^[��]ËL$�A   �   t2�D$�H�3��f��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�d�5    �B	3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�u�Q�R9Qu�   �SQ�0U	�SQ�0U	�L$�K�C�kUQPXY]Y[� �������������������������������������������������������������������������������̋�U���S�u�M��hM���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�
?��YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�vP���� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�����������������������������������������������̋�U��=�o	 u�E��N	�A#E]�j �u�u��Y����]������������̋�U��UV�u�23�;�r;�s3�@�U�
^]���������̋�U��E�jY#�U����  �yJ���B+ʃ����M�҅�t
3�]Ã<� u�@��|�3�@]������������������̋�U��ESVW�jY#�U����  �yJ���B�}+�3�B���3ۍ4;�r;�s3�C�4����t���Q3�;�r��s3�C��Hy�_^��[]���������������������������̋�U��QQ�e� SVW�}O�G�����G��%  �yH���@�ujY+�3�@���M�����   �������҅���<� u@��|��e�ǙjY#������  �yO���G�e 3�+�B����<;�r;�s�E   �M�<����t���Q3�;�r��s3�G����Hy��M��M������jY!�C;�}	+ˍ<�3��E�_^[������������������������������������������������������������̋�U��E�MjZ+�V�0�4��Ju�^]�������̋�U��W�}3����_]����̋�U��3��M�<� u@��|�3�@]�3�]�������̋�U��E�����UV����  �WyJ���B�e� �e �}��������E�    )U�S�֋M��#މ]������M]����]�M����E�}�]�|�jY��+Ѝ�[;�|�2�4���$� ��Iy�_^���������������������������������������̋�U���<�B	3ŉE��E�M�M��H
�с� �  �MċH�M��H� S�]���  ���?  ��VW�U��M�E������u"3�3�9t��u@��|��  3��}𫫫�3  �e� �u��}䥥�¥�{�E�O�G�������W��  ��E�yJ���B�t��j3�Y+�@���M̅��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}܋99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U܉�M�yщMЋM̃����jY!�E�@;�}
�|��+�3��}� t�E��C�M���+S;�}3��}𫫫�  ;��  +Eԍu�}𥥋ș����4������  �yJ���B�e� �e� ��������E�    )U��ЋM��|����#ȉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���E�Y+�;�|��T����d�� ��Iy�{O�G�������W��  ��E�yJ���BjY+�3�B��M̅T����   �������օt����|�� uB��|��o�ǙjY#������  �yO���G�e� 3�+�B��L���9�4�u�;�r;�s�E�   �U܉�M����t�L����r3�;�r��s3�G�1��HyދEԋM̃����jY!T��@;�}
�|��+�3��K�A����4�Q����  �yJ���B�e� �e� ��������E�    )U��ЋM��|����#ȉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���E�Y+�;�|��T����d�� ��Iy�3�jX�N  ;�K��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�s33�@�   �su��e�������������с�  ��E�yJ���B�e� �e� ��������E�    )U��׋E��D����#ωMԋ���M�E؉D���EԋM����E��}��E�|ЋŰ�j���E�Y+�;�|�8�|����d�� ��Iy�3�jY+K�[��M���Ɂ�   ��u���@u�MȋU�q��
�� u�Mȉ1�M�_^3�[�[������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�B	3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=LU	O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�HU	��+LU	;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5LU	N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��PU	�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �PU	;DU	��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�XU	DU	3�@�   XU	�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+PU	��M���Ɂ�   �ًTU	]���@u�M̋U�Y��
�� u�M̉�M�_3�[��T�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���8�B	3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=dU	O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�`U	��+dU	;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5dU	N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��hU	�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �hU	;\U	��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�pU	\U	3�@�   pU	�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+hU	��M���Ɂ�   �ًlU	]���@u�M̋U�Y��
�� u�M̉�M�_3�[�JN�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��� �B	3ŉE��M�Q
�e� ��%�  �� �  V�q�E�Q�	��W�}�u��M���yd�����t\�J3�;�r��s3�F�e� �M�΅�t8�M�e� �L����r;�r��s�E�   �M�1�M�y҅�t
�E�   ���u��U���  f9M�u�E�   E�M��wf�G�E��_3�^�L����������������������������������������������������������̋�U��EV�0���W�x���0�4?�H������_�p�H^]������������̋�U��E�P�HVW��������ΉH��������_�P�^]������������̋�U���0�B	3ŉE��E3�S�]�S
V�MԉM��M�M��H
��3�� �  �u��  #�#֍4
W����  �u�f;���  f;���  ���  f;���  ��?  f;�w
3ɉH��  ����f��uF�uЅxu3�9Hu9uf�H
�  3�f;�uF�uЅ{u	9Ku9t��M�}��E�   �M�U�ɉU؅�~P���]܍�U����e� �ʋW��4
;�r;�s�E�   �}� �w�tf��m����M؃}� ��]�uЃ��E��M�}� ����  ���  f��~8�E�   �u*�M��]�U��e����ًM�������]�M�f���f��O�f��yH�����ɉM���E�t�EԋM��]�U��m�����ًM�������M�]�M�uσ}� tf�M�� �  f9M�w�U����� �� � u/�}��u&�e� �}��u�e� f9}�uf�M�F�f�E���E���E��  f;�sf�M�u�f��M�H�M��Hf�p
� 3�3�f9M���J��   ��� ���P��H�M�_^3�[��H�����������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���D�B	3ŉE��E��U	��`3҉M�9U��  }�]��V	��`�M�9Uu3�f�9U��  SVW�M�E�T�}��;��~  k�M܋ٹ �  f9r��}䥥��M�]��H
�UȉU��U�U��S
��3�� �  �uо�  #�#֍<
���}�f;��  f;���  ���  f;���  ��?  f;�w
3ɉH��  3�f;�u!G�@����}�u9pu90u3�f�H
��  f;�u#G�C����}�u9su93u�p�p�0�  �u̍u��E�   �M̋U�ɉUԅ�~S�SȉU��MċMċU���	�e� �ʋV��<
;�r;�s�E�   �}� �~�tf��E��m��Mԃ}� ��}؃��E��M��}� ����  f��~;�E�   �u-�u�M��e�������M����ʁ���  �u�M�f���f��M����  f��yB��������E�t�EȋM��]�U��m�����ًM������N�]�M�u�9u�tf�M�� �  f9M�w�U����� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�M�G�f�E���E���E��  f;�sf�M�}�f��M�H�M��Hf�x
� 3�3�f9M���J��   ��� ���P�H�3�9U�a���_^[�M�3��ME��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���|�B	3ŉE��E3�V3��E��EFW�E��}��M��u��M��M��M��M��M��M��M�9M$u�W@���    ��@��3��<  �U�U��< t<	t<
t<uB��S�0�B���  �$���Hπ�wjYJ�ߋM$�	���   �	:ujY������+tHHt���|  ���jY�E� �  뤃e� jY뛍Hωu���v��M$�	���   �	:uj�<+t"<-t:�t�<C�/  <E~
,d<�!  j�Jj넍Hπ��_����M$�	���   �	:�a���:��s����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�h���<+t�<-t��k����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Hπ�wj	��������+t HHt���=���j�����M��jY�Q���j�~����u���B:�t�,1<v�J�&�Hπ�v�:�뿃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�]����B:�}��Q����M��E�O�? t�E�P�u��E�P�^#���E�3҃�9U�}��E�9U�uE9U�u+E=P  �!  =�����-  ��U	��`�E�;���  }�ع�V	�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k��� �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��   f;��  ���  f;��	  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� ����E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��yB��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  f9E�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �=����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W[�M�_3�^��=���ÍI ҭ$�o�����1���u�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����B	3ŉE��U�M�EV�uWR3�RRR�uQP�E�P�.�����E�VP�)����(��u���M���_3�^�;�������������������������̋�U��E�SVW�}��43�;�r;�s3�C�0��t�H�Q3�;�r��s3�F�P��t�@�H�W�43�;�r;�s3�C�p��t�@�OH_^[]����������������������������̋�U���t�B	3ŉE��E�U� �  #�S�]�E��A�V#�f�}� W�]��E������E������E����?�E�   t�C-��C �u�}f��u7����   ����   3�f9M�f�����$ �Cf�C0�C 3�@�  f;���   �M3�@f��   �;�u�} t��   @uh�	�S3�PPPPP��,��3�f9U�t��   �u9Uu-h�	�;�u"9Uuh�	�CjP�s7������u��C�h�	�CjP�V7������u��C3��k  �ʋ�i�M  �������Ck�M��������3�f�M��ع�U	��`�ۉE�f�U�u�}�M���  ��y��V	��`�ۉE�����  �E�T�������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E����E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��yB��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��}����M�����?  ��  f;���  �]��E�3҉U��U��U�U��U�3�#�#Ё� �  �4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��Z���3�3�f9u���H%   � ���E��a���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~K�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m����M��}� ����E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��yB��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t0����)3�f�� �  f9E�f�B0����$ �B�B �s�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�y2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K����C���<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[�B2���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��QQ�EV3��} 	 u:���u5��}��M���=  �=  f;�u95��	t5�]��M�����  ���  t %����P�uV�� ������t
VVVVV�5"��^�����������������������������̋�U��M3���tjX��t����t����t���� t����t   S��V�ʾ   #�W�   �   t!��   t��   t;�u��	��   #�t;�u   �   �E   _^[t   ]����������������������������������������3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �����������������������������������̋�U��M3���?t2��tjX��t����t����t���� t����t   ]�����������������3���yjXS�   VW��t����   t����   t����   t���   ��t   �ʾ `  #�t!��    t�� @  t;�u   ����_��@�  ��@^[t���  t��@u   �   �   �����������������������������������������3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  ����������������������������������������̋�U��M3���?t2��tjX��t����t����t���� t����t   ]�����������������h�  �T��Y���̋�U��QQV��}��E�3Ҿ   �?t)�tjZ�t���t���t��� t���tփ=��	 tA�]��M�3���?t/��tjX��t����t����t���� t����t�����^�������������������������������������̋�V�����0���5���h�  �~ ��Y��t�F�   t�`  �@$��  ^������������������3ɨ?t-�tjY�t���t���t��� t���t��   ����������������̋�U��Q�]��e���U��M�3���?t2��tjX��t����t����t���� t����t   ���������������������̋�U��QQ�e�]��M�3���yjXS�   VW��t����   t����   t����   t���   ��t   �ѿ `  #�t!��    t�� @  t;�u   ���ƾ@�  #΃�@t���  t��@u   �   �   �U�M#M��#��;���   �]���P�E������Y�]��U�3���yjX��t����   t����   t����   t���   ��t   ��#�t$��    t�� @  t;�u   �	   ��#փ�@t���  t��@u   �   �   _^[����������������������������������������������������������������������������������������������̋�U��U��t<��}�E3ɨ?t-�tjY�t���t���t��� t���t��   �
V�u��t�+����^]����������������������̋�U��QQ�}���=��	 ��   �E�3�V�   �?t)�tjZ�t���t���t��� t���t��]��e���U��M�3���?t/��tjX��t����t����t���� t����t��^�ÊM�3���?t2��tjX��t����t����t���� t����t   �������������������������������������������������������̋�U��E��SV3�W�   9U�V  ��}�f�]���tjZ��t����t����t���� t����t��   �ËȾ   #�t&��   t��   t;�u����   ���   #�t=   u��   ���   �é   t��   �]�E#E��#��;���   �=������E��m���}��U�3���tj[��t����t����t���� t����t��   �ʋ�#�t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �E��E�} ��  3�95��	�~  %�E��]�E��yj^�   t���   t���   t���   t���   t��   �ȿ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #Ã�@t-�  t��@u��   ���   ���   �E���#E��#��;�u���   ����P�E�����Y�]�M3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#˃�@t���  t��@u��   ���   ���   �M���E�0_3�^@[������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���SVW��}�f�]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   �é   t��   �}�M����#�#���E;���   ���h������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95��	��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��"���Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U���SVW�}��������}f�]3���tjZ��t����t����t���� t����t��   �ˋ��   #�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   �é   t��   ���Ћ�#M#���E�;���   ���������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U�3�95��	��  ���}��]�E��yj^�   t���   t���   t���   t���   t��   �ȿ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #Ã�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   �����P�E��C���Y�]��U�3���yjX��   t����   t����   t����   t���   ��t   ��#�t$��    t�� @  t;�u   �	   ��#Ӄ�@t���  t��@u   �   �   ��3M�E��� t   �_^[������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��EVW��xY;T�	sQ���������<���	����<�u5�=`_	S�]u�� tHtHuSj��Sj��Sj��ܒ	��3�[����� 	   �h����  ���_^]��������������������������������̋�U��MS3�VW;�|[;T�	sS��������<���	����D0t6�<0�t0�=`_	u+�tItIuSj��Sj��Sj��ܒ	���3������� 	   ���������_^[]���������������������������������̋�U��E���u�����  ���� 	   ���]Å�x;T�	r�a����  ���� 	   �)���Ջ�������	�����Dt͋]���������������������������jh�,	�	���}����������4���	�E�   3�9^u5j
����Y�]�9^uh�  �FP�4�	��u�]��F�E������0   9]�t������������	�D8P���	�E��G���3ۋ}j
���Y���������������������������������������̋�U��E�ȃ�������	���DP���	]����������jh�,	����M��3��}�j�!���Y��u����a  j����Y�}��}؃�@�;  �4���	����   �u�����	   ;���   �Fu[�~ u8j
�]���Y3�C�]��~ uh�  �FP�4�	��u�]���F�e� �(   �}� u�^S���	�FtS���	��@냋}؋u�j
����YÃ}� u��F��+4���	��������u�}��uyG�,���j@j �s��YY�E���ta����	��T�	 ���   ;�s�@ ���@
�` ��@�E������}�����σ�������	�DW�R���Y��u�M���E������	   �E��R���j���Y�������������������������������������������������������������������������������������������������������jh(-	���3��}�2��Et�� �E @  t�ˀ�E�t���u�8�	;�u��	P����Y������Ã�u��@���u���$�����u���u�����    �����8�}��uV���YY����������	�ƃ�����\��T$�"��	�D$� �E�   �E������   9}��i������e����u3�9}�u�����΃�������	�D� �V����Y���������������������������������������������������������������������̋�U��Q�=�X	�u������X	���u���  ��j �M�Qj�MQP���	��t�f�E������������������jhH-	�b��j����Y�e� �u���Y���E��E������
   f�E��� ���j���Y�����������������̋�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M������E�9Xu�E;�t�f�8]�t�E��`p�3�@�ˍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�Ԓ	���E�u�M;��   r 8^t���   8]��f����M��ap��Z����r��� *   8]�t�E��`p�����;���3�9]��P�u�E�jVj	�p�Ԓ	���:������������������������������������������������������������������������̋�U��j �u�u�u�z����]�������jhh-	���3ۉ]�j�@���Y�]�j_�}�;= �	}T����o	9�tE���@�tP�����Y���t�E��|(��o	���� P�@�	��o	�4����Y��o	��G��E������	   �E�������j����Y���������������������������������������̋�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV����YP������;�u�F��y����F��N ���_�F�f �^��[]��������������������������̋�U��V�u��u	V�G   Y�/V�-
��Y��t�����F @  tV�+���P�����Y��Y��3�^]�������������������jh�-	�� ��3��}�}�j����Y�}�3��u�;5 �	��   ��o	��98t^� �@�tVPV���YY3�B�U���o	���H���t/9UuP����Y���t�E��9}u��tP���Y���u	E܉}��   F�3��u��o	�4�V���YY��E������   �}�E�t�E�������j����Y�������������������������������������������������������jh�-	�����3�9uu	V�����Y�'�u�����Y�u��u� ��Y�E��E������	   �E��l�����u�Y��Y���������������������j����Y��̋�U��V�uV�u���P���YY��t|�<����� ;�u3���,�����@;�u`3�@��o	�F  uNSW�<��o	�? �   u S�����Y���u�Fj�F�X�F�F��?�~�>�^�^�N  3�_@[�3�^]���������������������������������������̋�U��} t'V�u�F   tV����f�����f �& �f Y^]��������������jh�-	�k����G����p �u�3�9E����u�
���    �#������<V�X���Y�e� V�������u�u�uV�U�E�VW������E������   �E������Ëu�V����Y���������������������������������̋�U���u�u�uh��������]�������̋�U���u�u�uh���������]�������̋�U���u�u�uh�������]�������̋�U���uj �uh��������]�������̋�U���uj �uh���t�����]�������̋�U���uj �uh��Q�����]�������̋�U���V�u�M��"����E�u��t�0��u$�	���    �	���}� t�E�`p�3���  �} t�}|Ѓ}$ʃe� �M�S�W�~���   ~�E�P��jP����M������   ���B����t�G�ǀ�-u�M���+u�G�E���O  ���F  ��$�=  ��u*��0t	�E
   �6�<xt<Xt	�E   �#�E   �
��u��0u�<xt<Xu�_�����3��u���   �U����N�у�t�˃�0���  t0�K�����w�� ���;Ms�M9E�r(u;M�v!�M�} u#�EO�u �} t�}�e� �[�U��UщU��G늾����u�u=��t	�}�   �w	��u+9u�v&�c���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�_[^�������������������������������������������������������������������������������������������������������������������������������������������̋�U��3�P�u�u�u9�o	uh�N	�P�%�����]����������̋�U��j �u�u�u�u�������]�������̋�U��=�o	 j�u�u�uuh�N	�j �������]�����������̋�U��j�u�u�u�u������]�������̋�U���<S�u�M������M�E3�;�t�;�u%����    �<��8]�t�Ẽ`p�3�3��O  9]t�}|Ѓ}$ʊV�u�W�]�]��M��x���   ~�E�P�E�jP�����uă���E����   �A��;�t��E�G�}�-�}�u�M��}�+u	�G�}��E�jY9]u%�}�0t	�E
   �7�<xt<Xt	�E   �$�M9Mu�}�0u�<xt<Xu�G���E��}��E�R��Wj�j��U������]����   �M܉E�U�M����C�Ѓ�t���0�%  tP�A�<��w�� �p�;us;�M��M;M�rQw�E�;E�rG�E�9E�u;M�u3�;E�r3w;u�v,�M�} u;�E�M��uA3�9Et�M�M��E�E��   Q�u��u�W�.���3��щE�U��E�� �E��E��E��������   ��u'�uT��t9]�wr�}� w��u>9u�r9w�}��v1����E� "   t
�M���M����Et	�e� �]���M���u��E_^��t�M���Et�E�M��؃� �ىE�M��}� t�Ẽ`p��E�U�[������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��3�P�u�u�u9�o	uh�N	�P������]����������̋�U��j �u�u�u�u�o�����]�������̋�U��=�o	 j�u�u�uuh�N	�j �<�����]�����������̋�U��j�u�u�u�u������]�������̋�U���S�u�M�������M3�;�u8]�t�E��`p�3��   9]u&����    �5��8]�t�E��`p������   9]t�V����;�v�\���    � ���?�E�9Xu�uQ�u�u��������6�pQ�uQ�uh  �p�E�P�>����� ;�u8]�t�E��`p�������8]�t�M��ap�^[��������������������������������������������������������̋�U��j �u�u�u������]������̋�U��QQSV3�W�=�_	�u��;�te�L�	VVVVj�PVV�ӉE�;�tTjP���YY�E�;�tCVV�u�Pj��7VV�Ӆ�t6�E�VP���YY��y9u�t�u������Y�u����;�u�3�_^[�Ã�����u������Y��������������������������������������̋�U��Q�e� V�E�P�u�u����������u9E�t������t
�����M����^�����������������̋�U��3�9Ev�M�9 t@A;Er�]��������3�Ë�U��MVW��t�}��u�I���j^�0��������A�U��u� ���> tFOu���t�+��B��tOu��u� ����j"Y����3�_^]���������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������������̋�U��3�S3�@9]|FVW��t>�EÙ+��E���<��7�E�0�����YY��u
�M���9�yN�u��^;]~�_^3Ʌ���[��]������������������������́N  ��	�F�F�����̋�U��Q��tP�> tKh	V�����YY��t:h	V����YY��uj�E�Ph   �w���	��t)�E���V�����Y�E���j�E�Ph  �w���	��u3��Ã}� u����	����������������������������������̋�U��3�f�Mf;��	t����r�3�@]�3�]���������̋�V3�� �A�B<w����
�A�<w�������t�Њ
��uڋ�^�������������3��
B��A|��Z~��a��w@��������̋�U���|�B	3ŉE�VW�}�����׋��}�����jx�E�P���   ���%���  PW��	��u	!��   @�A�E�P���   ����YY��uW����Y��t���   ���   ���   ���   ���Ѓ��M�_3�^�  ���� ����������������������������������������̋�U��QV��j�E�P��%�  h      P���	��u3��);u�t!�} t�E�0W�������V���*���Y;�_t�3�@^�����������������������̋�U���|�B	3ŉE�SVW�}������׍��   �7�����	��jx�E�P�F���%���  PW�Ӆ�u�f 3�@�c  �E�P�v����YY����   jx�E�P�F���%���  PW�Ӆ�t��E�P�6����YY��u�N  �~�R�FuO�F��t,P�E�P�6�e�������u�6�N�~�+���Y;Fu!�~��V��uW�=���Y��t	���V�~�N�   #�;���   jx�E�P�F���%���  PW�Ӆ������E�P�6�����Y3�Y��u0�N   �F9^t
   �F�H9^t<�6����Y;Fu/Vj�9^u49^t/�E�P�6����YY��uVS�������YY��t�N   9^u�~�F���Ѓ��M�_^3�[������ �������������������������������������������������������������������������������������������������������������������̋�U���|�B	3ŉE�VW�}�����׍��   �������jx�E�P�F���%���  PW��	��u!F@�\�E�P�6����YY��u
9Fu1Vj��~ u0�~ t*�E�P�6�Z���YY��uVP������YY��t
�N�~�~�F���Ѓ��M�_3�^�a����� �������������������������������������������������v���������Y�j@h+��F��	�Fu�f �������������6�����v�����@�F����������f @�~ YY�FtjX�������jhl��F��	�F�   t�   t�u�f ���������������������������6���������@Y�FtjX������jh���F��	�Fu�f ���������������̋�U��SVW�������   �E��u�O  ��   ���@�_�t�8 tSjh 	��������g ��t[�8 tV���t�8 t	�����������D���� ��   Wj@h�	�<�������tf���t�; t	�������R�������I���t0�; t+S��������Y�j@h+��G��	�Gu�g ��G  ��	�G�G� ��   �u�ƃ����#��E������u����   ����  ��   ����  ��   ��P���	����   j�w��	����   �E��tf�Of�f�Of�Hf�p�]��th�5�	�  f9u h	j@S��������t3�PPPPP�^���j@Sh  �w�օ�t,j@�C@Ph  �w�օ�tj
j��S�u������3�@�3�_^[]����������������������������������������������������������������������������������������������������������������������������̅�t3Ʌ����D	������� �	+�t3Ʌ����D	�������f�f;t1���+�t3҅��D���u�F�I+�t3Ʌ����D	��3����������������̋;tg���+�t3҅��D���uP�F�Q+�t3҅��D���u5�F�Q+�t3҅��D���u�F�I+�t3Ʌ����D	��3�����������������������������̋�VW���N  �;tv���+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������t ����3�����  �A;Btw���B+�t3������D ����k  �q�B+�t3������D ����L  �q�B+�t3������D ����-  �q�B+�t3������t ����3����  �A;Btw���B+�t3������D �����  �q	�B	+�t3������D �����  �q
�B
+�t3������D �����  �q�B+�t3������t ����3����  �A;Btw���B+�t3������D ����Y  �q�B+�t3������D ����:  �q�B+�t3������D ����  �q�B+�t3������t ����3�����  �A;Btw���B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������t ����3����m  �A;Btw���B+�t3������D ����G  �q�B+�t3������D ����(  �q�B+�t3������D ����	  �q�B+�t3������t ����3�����  �A;Btw���B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������D �����  �q�B+�t3������t ����3����[  �A;Btw���B+�t3������D ����5  �q�B+�t3������D ����  �q�B+�t3������D �����  �q�B+�t3������t ����3�����  �� �� �� �� ������׃���  �$���A�;B�tx�B��q�+�t3������D �����  �q��B�+�t3������D ����f  �q��B�+�t3������D ����G  �q��B�+�t3������t ����3����"  �A�;B�tw���B�+�t3������D �����  �q��B�+�t3������D �����  �q��B�+�t3������D �����  �q��B�+�t3������t ����3�����  �A�;B�tw���B�+�t3������D ����s  �q��B�+�t3������D ����T  �q��B�+�t3������D ����5  �q��B�+�t3������t ����3����  �A�;B�tw���B�+�t3������D �����  �q��B�+�t3������D �����  �q��B�+�t3������D �����  �q��B�+�t3������t ����3�����  �A�;B�tw���B�+�t3������D ����a  �q��B�+�t3������D ����B  �q��B�+�t3������D ����#  �q��B�+�t3������t ����3�����   �A�;B�tw���B�+�t3������D �����   �q��B�+�t3������D �����   �q��B�+�t3������D �����   �q��B�+�t3������t ����3���uy�A�;B�ti���B�+�t3������D ���uW�q��B�+�t3������D ���u<�q��B�+�t3������D ���u!�A��J�+�t3Ʌ����D	��3���u3�_^ËA�;B�tk���B�+�t3������D ���u��q��B�+�t3������D ���u��q��B�+�t3������D ���u��q��B�+�t3������t ����3���u��A�;B�tx�B��q�+�t3������D ����]����q��B�+�t3������D ����>����q��B�+�t3������D ��������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3����q����A�;B�tw���B�+�t3������D ����K����q��B�+�t3������D ����,����q��B�+�t3������D ��������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3����_����A�;B�tw���B�+�t3������D ����9����q��B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ����r����q��B�+�t3������t ����3����M����A��J�+��=���3Ʌ����D	��-����A�;B�tw���B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tx�B��q�+�t3������D ����}����q��B�+�t3������D ����^����q��B�+�t3������D ����?����q��B�+�t3������t ����3��������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ����k����q��B�+�t3������D ����L����q��B�+�t3������D ����-����q��B�+�t3������t ����3��������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3��������A�;B�tw���B�+�t3������D ����Y����q��B�+�t3������D ����:����q��B�+�t3������D ��������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3����m���f�A�f;B��]�����  �A�;B�tx�B��q�+�t3������D ����3����q��B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ����l����q��B�+�t3������t ����3����G����A�;B�tw���B�+�t3������D ����!����q��B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ����y����q��B�+�t3������D ����Z����q��B�+�t3������t ����3����5����A�;B�tw���B�+�t3������D ��������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3���������A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ����g����q��B�+�t3������D ����H����q��B�+�t3������t ����3����#����A�;B�tw���B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������D ���������q��B�+�t3������t ����3���������q��B�+�t3������D ����{����q��B�+�����3������D ������6��	��bB	:���� P0( ��z��>�
���h
��;�	�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��VW�}�ǃ� ��  H��  H�l  H�!  H��  �M�ESj Z�2  �0;1tt�0�+�t3ۅ��Ít����+  �p�Y+�t3ۅ��Ít����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����e  �p�Y+�t3ۅ��Ít��3����B  �p;qtv�p�Y+�t3ۅ��Ít����  �p	�Y	+�t3ۅ��Ít�����  �p
�Y
+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����t  �p�Y+�t3ۅ��Ít����U  �p�Y+�t3ۅ��Ít��3����2  �p;qtv�Y�p+�t3ۅ��Ít����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����d  �p�Y+�t3ۅ��Ít����E  �p�Y+�t3ۅ��Ít��3����"  �p;qtv�p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít��3�����   �p;qtj�p�Y+�t3ۅ��Ít���uw�p�Y+�t3ۅ��Ít���u\�p�Y+�t3ۅ��Ít���uA�p�Y+�t3ۅ��Ít��3���u"��+�;�������σ���  �$�D(���  �P�;Q�ti���Q�+�t3҅��t���u��p��Q�+�t3҅��t���u��p��Q�+�t3҅��t���u��p��Q�+�t3҅��t��3���u��P�;Q�tu���Q�+�t3҅��t����\����p��Q�+�t3҅��t����=����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����t����P�;Q�tu���Q�+�t3҅��t����N����p��Q�+�t3҅��t����/����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����e����P�;Q�tu���Q�+�t3҅��t����?����p��Q�+�t3҅��t���� ����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tm���Q�+�t3҅��T���u6�p��Q�+�t3҅��T���u�p��Q�+�t3҅��T���t����@��I�+�t3Ʌ����D	��3���u3�[�  �P�;Q�tu���Q�+�t3҅��t����5����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t����p����p��Q�+�t3҅��t��3����M����P�;Q�tu���Q�+�t3҅��t����'����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t����b����p��Q�+�t3҅��t��3����?����P�;Q�tu���Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������p��Q�+�t3҅��t����r����p��Q�+�t3҅��t����S����p��Q�+�t3҅��t��3����0����P�;Q�tu���Q�+�t3҅��t����
����p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������I��@�+��8���3Ʌ����D	��(����P�;Q�tu���Q�+�t3҅��t����c����p��Q�+�t3҅��t����D����p��Q�+�t3҅��t����%����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����{����P�;Q�tu���Q�+�t3҅��t����U����p��Q�+�t3҅��t����6����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����m����P�;Q�tu���Q�+�t3҅��t����G����p��Q�+�t3҅��t����(����p��Q�+�t3҅��t����	����p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������Q��p�+�t3҅��t���������Q��p�+�t3҅��t���������Q��p�+�t3҅��t��3����^����P�;Q�tu���Q�+�t3҅��t����8����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3��������f�P�f;Q��f����Q��p�+�����3҅��T�����  ������P�;Q�tv�Q��p�+�t3҅��t����z����p��Q�+�t3҅��t����[����p��Q�+�t3҅��t����<����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t����l����p��Q�+�t3҅��t����M����p��Q�+�t3҅��t����.����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t����]����p��Q�+�t3҅��t����>����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����u����P�;Q�tu���Q�+�t3҅��t����O����p��Q�+�t3҅��t����0����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������p��Q�+�����3҅��T����������c����M�u��+�t3҅��D�����   �A�V+�t3҅��D�����   �A�V+�t3҅��D�����   �A�N+���   3Ʌ����D	��   �M�u��+�t3҅��D���ud�A�V+�t3҅��D���uI�A�N뤋M�u��+�t3҅��D���u �A�N�x����E�M� �	�g���3�_^]Ë��U'#' ��"�&�F"&��!z%�8
!�$�� l$|*��#�u]#��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��Q�e� S�]��u3��   V��ru�s���tn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9u�r��.�@��I��F�@��I��<�@��I��2�@��I��(�M�E�u�����t:u@FA;�r�3�^[��� �	+����������������������������������������������������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�����������������̋�U����ES3�VW�E�N@  ��X�X9]�E  �]����}襥��э<	���ʋU�e ��ى}����֋u����ϋ��M���U�����։0�x�H;�r;U�s�E   �} �t'�u��e �~;�r��s�E   �} �xtA�H�u�e �7;�r;�s�E   �} �XtA�HM��e� ��ɋ��������މH�M�M�M��X�1�2�u�;�r;�s�E�   �}� �t$�K3�;�r��s3�B�ىH��t
�M�A�M�H�M�M�E�} �X�H�����3�9Xu*�P��E���  ��������������P�;�t܉x�x�� �  u0�H��E���  �����������ʉ�H�x�� �  t�f�M�_^f�H
[���������������������������������������������������������������������������������������������������������������������������3�PPjPjh   @h4	���	��X	�������̡�X	���t���tP���	�����̋�U��V�uW�����u�ѻ���    �u�����D�F�t8V�x���V���U���V聦��P��������y�����F��tP�N����f Y�f ��_^]����������������������������jh�-	�#����M��3��u������u�<����    ���������F@t�f �E�豫���V����Y�e� V�x���Y�E��E������   �ԋuV�z���Y������������������������������jh.	蒮���]���u赺��� 	   ����   ��x;T�	r薺��� 	   �:����ڋ����<���	�������D��t�S�ݐ��Y�e� ��Dt1S�|���YP���	��u��	�E���e� �}� t������M������ 	   �M���E������   �E�蘪��Ë]S�{���Y��������������������������������������������������������A@t�y t$�Ix��������QP�y���YY���u	��������������̋�U��V����M�E�M�����>�t�} �^]���������̋�U��QSV�����@����G@� �E�t
� u�J�&����  �(�E� ��K�U����E�>�u�����8*u�ϰ?�:�����������8 u
�����M��^[������������������������������̋�U���x  �B	3ŉE�S�]V�u3�W�u�}�������������������������������������������������������������c�����u+�P����    ����������� t
�������`p�����	  �F@u^V�����Y�`B	���t���t�ȃ����������	����A$u����t���t�ȃ��������	����@$��q���3�;��g�������������������������������������Z
  G������9������1
  �B�<Xw����(	���3�������k�	��H	j��^������;������jY;���	  �$��@3���������������������������������������������	  �� tH��t4+�t$HHt���q	  	������f	  �������Z	  �������N	  �������   �?	  �������3	  ��*u,���������[����������	  �������������	  ������k�
�ʍDЉ�������  ������ ��  ��*u&���������[�����������  ��������  ������k�
�ʍDЉ������  ��ItU��htD��lt��w�}  ������   �n  �?luG������   �������S  �������G  ������ �;  �<6u�4u�������� �  �������  <3u�2u�������������������  <d��  <i��  <o��  <u��  <x��  <X��  ������ ������ ������P��P�����Y��������Yt"�������������<����G������������������������������c  ��d��  �w  ��S��   ��   ��AtHHtYHHtHH��  �� ǅ����   ������������@������ �������   �������������E  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  �������[���������  ��u��E	������������ǅ����   �s  ��X��  HHty+��&���HH��  ��������  ������t0�C�Ph   ������P������P��������tǅ����   ��C�������ǅ����   �������������)  �����������t<�H��t5������   � ������t�+���ǅ����   ��  ������ ��  ��E	������P�r���Y��  ��p��  ��  ��e��  ��g�2�����itm��nt$��o��  �������������ta������   �U�3���������������"��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ދC��S���  u��gucǅ����   �W9�����~�������������   ~=��������]  V菆��������Y��������t���������������
ǅ�����   ��5ԑ	���������C�������������P��������������������P������������WP�58B	���Ћ���������   t������ u������PW�5DB	����YY������gu��u������PW�5@B	����YY�?-u������   G������W�����������������$��s�����HH���������  ǅ����'   �������ǅ����   �t���������Qƅ����0������ǅ����   �P�����   �V������� t��������@t�C���C����C���@t��3҉�������@t��|��s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW讘����0���������ڃ�9~������N뽍E�+�F������   ������������tc��t�΀90tX�������������0@�@If�8 t����u�+��������(��u��E	�������������I�8 t@��u�+����������������� �}  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+������������u'����~!������������� O������������t��ߋ�����������������P����������������Yt(������u��������ϰ0K�����������t��ヽ���� ������tT��~P�������Pj�E�P������PK���u�������u ��������t�E�P����������Y��u�������������������������t���Y������ |.������t%��������������ϰ K������������t��ヽ���� t�������>��������� Y���������������t������3������������� t����������������� t
�������`p��������M�_^3�[������Ë��8�6�6B7�7�7�79�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��S�]V�u�F<p�  ��p��   <st<St3��3�B��st	��St3��3�A����   ����   �d:�tM<it-<ot)<ut%<xt!<Xt:�t��it��ot��ut
��xt��Xu^:�t<it<ot<ut<xt<Xt3��3�A:�t��it��ot��ut��xt	��Xt3��3�@;�uK�F��3M��   u;3E� u4�3�;M���5;�u$�N�U�  #����#��������;�u3�@�3��	3�:�����^[]����������������������������������������������������������������������������A@t�y t$�Ix��������QP�A���YY���u	��������������̋�U��V����M�E�M�����>�t�} �^]���������̋�U��QSV���������G@� �E�t
� u�J�����  �(�E� ��K�U����E�>�u�ϧ���8*u�ϰ?�:������踧���8 u
讧���M��^[������������������������������̋�U��E� ��A��Q�]�����̋�U����  �B	3ŉE��ESV�uW�u�}3ۍ�������H�����������L�����������h�����D�����\����������������d���;�u*������    衧��8�����t
�������`p�����&  �F@u^V襑��Y�`B	���t���t�ȃ����������	����A$u����t���t�ȃ��������	����@$��r���;��j�����������4���������������u9������z  3ۋ�4�����l��������������������X�����`�����P�����p�������������������  ���������F������ ��|�����  �C�<Xw����(	���3���`���k�	��H	3���G3ɉ�`���;���   �>%��   �������uQj
��d���PV�x�������~2��d����8$u'������ uh@  ������j P�с����������������� 3�9�����u]j
��d���PV������d�����H������ �Q��������|���u(����  �9$��  ��d��  ;�l���~��l���3ɋ򋕀�����`����$�DY����  ���B  ��9�����u9������,  9������  ���������  �  ���������@�����D�����p�����h�����������\�����  �Ã� tI��t5��t%HHt����  �������  �������  	������  �������   �  �������  ��*��   9�����u�������������@��   j
��d���PV趄����d�����H������ �Q��|���uL����  �9$��  ������d�|  ;�l���~��l������Ŵ����9 ��   ������j*W�=  ���Ÿ���� 3ɉ�p���;���  ��������p����  ��p���k�
�ˍDЉ�p����  �������  ��*��   9�����u�������������@��<j
��d���PV�Ƀ����d�����H������ �Q��|����������Ÿ���� 3ɉ�����;��$  ��������  �9Ƅż���*���������������  ������k�
�ˍDЉ�������  ��ItU��htD��lt��w��  ������   �  �>luF������   ��|����  �������  ������ �  �<6u�~4u�������� �  ��|����c  <3u�~2u�������������|����A  <d��   <it|<otx<utt<xtp<Xtl��`�����\��� ������P��P�W��YY��t1��H������������������|���� ��|������������=  �؋�H����������������  ������   �  �Ã�d��  ��  ��S��   ��   ��AtHHtiHHtHH��	  �� ��@���������������@9�������  9�������  ��c��  �����Ŵ����9 �t  �   ��ż����	���������0  uw������   �k������0  u
������   ���������u����3�9������D  �������������@��}  ��X��  HH�&  ���7���HH��  ������  ��   9�����u�������������@��K��c��  9�����u.�����Ŵ����9 u�   ��  ������������j�)  ҋ�ո���� Ph   ������P��X���P��������tn��D����f9�����u�������������@��?��c�<  9�����u"�����Ŵ����9 u�9�V  �������  ҋ�ո���� ��������X����������������  9�����u�������������@�� ��c��  9�������   ҋ�ո���� ;�t8�H��t1������   � ������t�+�����\����N  ��\��� �B  ��E	������P��~��Y�+  ��p�   ��  ��e�  ��g�l�����i��   ��nt2��o��  ������ǅt���   ����   ��   �������   9�����u�������������p��C��c��   9�����u'�����Ŵ����9 ��  ������������j�>  ҋ�ո����0�!�������   ������ tf������f�����������D����>  ������@ǅt���
   ������3��� �  ��  9������D  ��������Q���������  ������������jQ����������  ������    裝�������� ����������� �������   ��������t���}ǅ����   �u4������gu������������ ud����������������@���8����o9�����~��������   9�����~���������]  V�q��Y��P�����t���������t�����듃�����c�-������������Ÿ������8����@�5ԑ	��<���������P��@���������������P��t�����8���SP�58B	���Ћ���������   t������ u������PS�5DB	����YY������gu��u������PS�5@B	����YY�;-u������   C������S����ǅ����   ǅL���   �$��s�����HH��������  ǅL���'   �������ǅt���   �������L���Qƅx���0��y���ǅh���   ������������c������9�����uu��Ŵ���91u�   �  S������j�L  ��   tZ9������k�����������c������9�����u$��Ŵ���91u�   �  S������j��   ��Ÿ�����Q�J  �� ��   ��@tJ9�����u�������������@���   ��������c�����9�������   ��Ÿ���� �   9�����u�������������@��   ��������c������9�����tD��Ÿ���� �n��@tl9�����u�������������@��O��������c������9�����u-��Ŵ���91��   S������WQ�]��������Z����*  ��Ÿ���� ��>9�����u�������������@��"��������c� ����9�����t���Ÿ���� 3���@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }'ǅ����   �5�9��������ż�����������~  ��������   9�����~���������u!�h��������������������������t-��t����RPSW�T�����0��X������ڃ�9~�L����N뽍�����+�F������   ��X�����������   ��t�΀90��   �������������0@��   ��c�����9�����u2�����Ŵ���91�����   ��������ż�����������   ҋ�ո���� ������  ������t4;�u��E	��������������\����	If90t��;�u�+��������,9�����u��E	�������������I�8 t@;�u�+�������X���������u������ ��  ��D��� ��  �������@t2�   t	ƅx���-��t	ƅx���+��tƅx��� ǅh���   ��p���+�X���+�h�����������t���u'����~!��H���������� O�����������t��ߋ�H�����h�����x���P�������Q���������Yt(������u��������ϰ0K�����������t��ヽ\��� ��X���tT��~P�������Pj�E�P��0���PK���r�������u ��0�����t�E�P�����������Y��u����������������������������Y������ |.������t%��t�����������ϰ K�����������t��ヽP��� t��P����;�����P��� Y��|�������������b���3�9�`���t��`����=���������uW9�����uO9�l���|G�������������H�ItItItItItItII������������F��������;�l���~�������������}3��q��������� t
�������`p��������M�_^3�[荘���Ð8IjI�I�I�J�J�K�L����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U��M�I�8 t@��u�I�E+�H]�������̋�U���,�B	3ŉE��ESVW�}�ىE܉U���~?��I�8 t@��u�������+���}�u��~*�΋�I�8 t@��u�������+���u����}�3���  ���|�e� �} u��@�E��t����   ;�ujX�  3�C;�~���  ;�~j��E�P�u���	��t���~-�}�r�}� �E�t؊P��tыM܊	:r:�v����8 u�뺅�~4�}�r��}� �E�t��P��t��M��	:r:��u������8 u��w����5Ԓ	j j W�u�j	�u�֋؉]ԅ������   ~@j�3�X���r4�D;�w�jq���ą�t� ��  �P�n��Y��t	� ��  ���E���e� �}� �����S�u��u�u�j�u�օ���   j j �u�u�j	�u�֋؅�tx~?j�3�X���r3�D;�w��p���ą�t� ��  �P�3n��Y��t	� ��  �����3���t1SW�u�u�j�u�օ�tSW�u��u��u�u� �	�E�W�<���Y�u��3����E�Y�e�_^[�M�3�����������������������������������������������������������������������������������������������������������������������������������������������������������������̋�U����u�M��x���u$�U�u �M��u�u�u�u��������}� t�M��ap������������������̋�U���S�u�M��=x���U3�;�u8]�t�E��`p�3��   9]u&�����    豌��8]�t�E��`p������   9]t�V����;�v�؋���    �|����K�E��H;�u�E�PR�u�u�\^�����?�p�E�R�uR�uh  QP�i���� ;�u膋���    8]�t�E��`p�������8]�t�M��ap�^[�����������������������������������������������������������̋�U��=�o	 u]��}��j �u�u�u�b����]����������̋�U��V�5�_	�!WP�u�:~������u��<=t��t�����uً�+�_	����^]Ë�+�_	�����������������������̋�U��QW��3��υ�tL9t	��@�9 u�V@jP蜌����YY�u���uj	�e���Y���t+�P��t������7Y��u�& �E�^_�������������������������̋�U����ES3ۉ]�;�u������    蜊������nV�0W�u�;�tSj=V�p����YY�}�;�t@;�t<3�8_���E���_	;�_	u
������_	;�u`9]t$9�_	t�]����tJ腉���    ���_^[��9]���  j�^��Y��_	;�tމ9�_	uj��]��Y��_	;�tÉ�5�_	�u�;�t�+}��u��8�����Y;�|R9tN�4��6�؇��Y9]�u�E���E��   �F��E�G�4�9u������?sjjW�5�_	�[����;�tU�N9]���   ;�}�ߍG;��6���=���?�+���Pj�5�_	�e[����;������U�����Y�M���_	9]tm�u�jV��h��Y��P蜊����YY;�tPVV��h��Y��PW躉������uR�M���+�E�@�����#�QW��	��u�M������� *   W�І��Y9]�t�u�����EY��E��s���SSSSS�~���u�袆���EY�3��T��������������������������������������������������������������������������������������������������������������������������������������������������̋�U����} SVW��   �u�M��*s���]��u'�����    踇���}� t�E��`p������   �u��tҿ���9}v!�܆���    耇���}� t�E��`p����]�E��x u�uVS�3[�����}� tA�M��ap��8+��3�M�QP�e������M�QP�e����F�Mt��t;�t�+����3�_^[���������������������������������������������������������̋�U��3�9�o	u09Eu�����    豆������]�9Et�}���w�]�mZ��P�u�u�u�X����]��������������������̋�U��SV��3�;�u諅��j^�0�P������   W9]w菅��j^�0�4������u3�9]���A9Mw	�l���j"�ۋM�����"wɋ�9]t3�C�-�N�؋�3��u��	v��W���0�AC��t;]r�;]r� �� I���I�G;�r�3�_^[]� ���������������������������������������������̋�U��}
�Eu
��yjj
�j �u�u�M�����]����������̋�U��3��}
u9E}@�MP�u�E�u����]���������̋�U��M�Ej �u�u����]������̋�U���3�V;�u�?���j^�0��������   9Mv�3�9M���@9Ew	����j"�ӋE�����"w��ES�]�M���9Mt����-�w�E�   �؉u�M�u�uPS��l���]��؋�	v��W���0��M�FA�M���u��t;MrȋM�[;Mr� 蒃��j"Y����L���� N�E���N�@�E;�r�3�^�� ����������������������������������������������������������̋�U��3��}
u9E
|9Es3�@W�}P�u�u�u�u����_]�������������̋�U��W�}j �u�u�u�u�{���_]�������̋�U��V�uWV��n��Y���tP���	��u	���   u��u�@Dtj�n��j���n��YY;�tV�n��YP���	��u
��	���3�V�ք����������	����Y�D0 ��tW��Z��Y����3�_^]����������������������������������������jh8.	��u���]���u�g���  ������ 	   ����   ��x;T�	r�g���  蹁��� 	   �]����ҋ����<���	�������D0��t�S� X��Y�e� ��D0tS�Ni��Y�E���g���� 	   �M���E������   �E���q��Ë]S��W��Y�������������������������������������������������̋�U��V�u�F��t�t�v����f����3�Y��F�F^]������������̋�U��S3�9]u3��>VW�u�Ba���pV�Ca����YY;�t�uVW��������u���SSSSS�Lw��3�_^[]��������������������̋�U���S�u�M��_l���E3�;�u �G����    ����8]�t�E��`p�3��pV�u�9^u:�uP�Ca��YY�=���D2t@�:�t:�������9MuH���9Ut	@�f;�u���9Mu8]�t�M��ap��8]�t�E��`p�3�^[���������������������������������������������̋�U��j �u�u�k����]�����������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��������������������������������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[������������������������������������������������������%̑	�%Б	�%ԑ	�%ؑ	�%ܑ	�%��	�%�	�%�	�%�	�%�	�%��	�%��	�%��	�% �	�%�	�%�	�%�	�%�	�%�	�%�	�%�	�% �	�%$�	�%(�	�%,�	�%0�	�%4�	�%8�	�%<�	�%@�	�%D�	�%H�	�%L�	�%P�	�%T�	�%X�	�%\�	�%`�	�%d�	�%h�	�%l�	�%p�	�%t�	�%x�	�%|�	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%��	�%Ē	�%Ȓ	�%̒	�%В	�%Ԓ	�%ؒ	�%ܒ	�%��	�%�	�%�	�%�	�%�	�%��	�%��	�%��	�% �	�%�	����U���@SVW�@Z	�ZQ��hЂ�W����_^[��]����������U���@SVWj �`Z	�*^��_^[��]���������������������U���@SVWh    jjj�z����P�z����P�	z������Z	_^[��]�����������������������U���@SVW��R����Z	_^[��]������̋�U��Q3��E���]����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������U���@SVW�@Z	��e��_^[��]�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �qr@r�r    �r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ������2�P�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                                                                                                                                                                                                                -�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ���P       o   �	 �T                                                                                                                                                                              	              	            	              	         ?             @                  �   &   ��������5            4  �������5            4  �������                                                 	       �������N���������������C-DT�!	@-DT�!�?        �������N���������������C-DT�!	@-DT�!�?        Ocontainer      Ocontainer.png          c:\program files\maxon\cinema 4d r14.025\plugins\_container object\src\containerobject.cpp                      d	��"�w�b�a�����%����������=�����T����H���������C����D��������                                ffffff�?              �?        333333�?             �o@                        �	��v�����f�������%����������=�����T����H���������C����D��������                                �	��v�����f�������%����������=�����                c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_resource.cpp                 #   M_EDITOR    �������N���������������C-DT�!	@-DT�!�?        res     �������N���������������C-DT�!	@-DT�!�?        �������?        -DT�!��              �        -DT�!�?              Y@        c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_memory.cpp                   �������N���������������C-DT�!	@-DT�!�?                c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_basebitmap.cpp               c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_misc\datastructures\basearray.h                      �������N���������������C-DT�!	@-DT�!�?        c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_file.cpp                     �������N���������������C-DT�!	@-DT�!�?        �	Y��� �e�����^� �(�        �������        ������             �f@        -DT�!	@             @�@     	���� �e�����^� ���        x 	�������K��������i�            c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_gui.cpp              � 	���� �e�����^� ���        ~       ,!	x��� �e�����^� ��z��������X�����y�	��                    Progress Thread     0%  %   �������N���������������C-DT�!	@-DT�!�?                ����MbP?    nncnt==ncnt     %s(%d): %s      nncnt<ncnt          c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_baseobject.cpp               �!	�{�    Stop    Stop:   c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_misc\datastructures\sort.h                   �!	�       %s      c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_general.h                    c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_pmain.cpp                    �������N���������������C-DT�!	@-DT�!�?              �?          4&�k�          4&�kC        c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_basetime.cpp                  �Ngm��C           ����A    �!	����]�]�        c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_libs\lib_ngon.cpp                    �������N���������������C-DT�!	@-DT�!�?        
   CRITICAL:       WARNING:     [%s %s L%d]    %H:%M:%S        c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_misc\memory\debugglobals.cpp                         c:\program files\maxon\cinema 4d r14.025\resource\_api\c4d_string.cpp               no baselist      B   KB  MB       �@     GB T"	��    ��                      �?      �?3      3            �      0C       �       ��                              fmod         ���;o;�;4;�;o;�;m;m;�;m;�;�;o;�;                                a/p am/pm   e+000   K E R N E L 3 2 . D L L         FlsFree     FlsSetValue     FlsGetValue     FlsAlloc    CorExitProcess      m s c o r e e . d l l         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �                                                                    �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ���5�h!����?      �?                            �?5�h!���>@�������             ��      �@      �                                          8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                r u n t i m e   e r r o r            
     T L O S S   e r r o r  
           S I N G   e r r o r  
         D O M A I N   e r r o r  
             R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
                                                                                                     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
                             R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
                                             R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
                     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
                 R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
                         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
                         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
                       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
                         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
                         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
                 R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
                         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
                           R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
                     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
                           R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
                       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
                            ��   x�	   �
   ��   @�   ��   ��   �   ��   8�   ��   8�   ��   ��   ��     �!   ��x   ��y   ��z   d��   \��   8�                                        M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y                 
 
     . . .       < p r o g r a m   n a m e   u n k n o w n >             R u n t i m e   E r r o r ! 
 
 P r o g r a m :                           �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��                    tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow �h	�h	    _nextafter      _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh        �������             ��      �@      �                    ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx                          H H : m m : s s         d d d d ,   M M M M   d d ,   y y y y           M M / d d / y y         P M     A M     D e c e m b e r         N o v e m b e r         O c t o b e r       S e p t e m b e r       A u g u s t     J u l y     J u n e     A p r i l       M a r c h       F e b r u a r y         J a n u a r y       D e c       N o v       O c t       S e p       A u g       J u l       J u n       M a y       A p r       M a r       F e b       J a n       S a t u r d a y         F r i d a y     T h u r s d a y         W e d n e s d a y       T u e s d a y       M o n d a y     S u n d a y     S a t       F r i       T h u       W e d       T u e       M o n       S u n       HH:mm:ss    dddd, MMMM dd, yyyy     MM/dd/yy    PM  AM  December    November    October     September   August  July    June    April   March   February    January     Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday     Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec                TZ   Complete Object Locator'        Class Hierarchy Descriptor'         Base Class Array'       Base Class Descriptor at (          Type Descriptor'       `local static thread guard'         `managed vector copy constructor iterator'          `vector vbase copy constructor iterator'            `vector copy constructor iterator'          `dynamic atexit destructor for '        `dynamic initializer for '      `eh vector vbase copy constructor iterator'         `eh vector copy constructor iterator'           `managed vector destructor iterator'        `managed vector constructor iterator'           `placement delete[] closure'        `placement delete closure'      `omni callsig'       delete[]    new[]  `local vftable constructor closure'         `local vftable'     `RTTI   `EH `udt returning'     `copy constructor closure'      `eh vector vbase constructor iterator'          `eh vector destructor iterator'         `eh vector constructor iterator'        `virtual displacement map'      `vector vbase constructor iterator'         `vector destructor iterator'        `vector constructor iterator'       `scalar deleting destructor'        `default constructor closure'       `vector deleting destructor'        `vbase destructor'      `string'    `local static guard'        `typeof'    `vcall'     `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete      new    __unaligned     __restrict      __ptr64     __eabi  __clrcall   __fastcall      __thiscall      __stdcall   __pascal    __cdecl     __based(        ����������������t�d�T�R�L�@�<�8�4�0�,�(�$������� �������\�������������е����������������������������������t�X�L�4����������T�4����������|�t�`�4�,� ��������l�<��������`�,��R���������p�                                                                                ]�]�]�    ������    }�����    :�����    ��H���    ����?�     ??     {flat}  {for    `non-type-template-parameter        unsigned    long    int     short   char    void    <ellipsis>      ... ,<ellipsis>     ,...     throw(     )[  s   '   `template-parameter     NULL    cli::pin_ptr<   cli::array<     void    ''  `anonymous namespace'       `   generic-type-   template-parameter-     ::  `unknown ecsu'      union   struct      class   enum    coclass     cointerface     )   extern "C"      [thunk]:    public:     protected:      private:    virtual     static      `template static data member destructor helper'             `template static data member constructor helper'            `local static destructor helper'        `adjustor{      `vtordisp{      `vtordispex{        }'  }'  const   volatile    CV:     volatile     volatile   const   signed      double  bool    <unknown>   wchar_t     UNKNOWN     __int128    __int32     __int64     __int16     __w64   __int8  float   long    int short   char    std::nullptr_t      SystemFunction036       A D V A P I 3 2 . D L L         GetProcessWindowStation     GetUserObjectInformationW       GetLastActivePopup      GetActiveWindow     MessageBoxW     U S E R 3 2 . D L L                                                                                                                                                                                                                                                                                           ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                            LC_TIME     LC_NUMERIC      LC_MONETARY     LC_CTYPE    LC_COLLATE      LC_ALL      �	    ���	L	���	L	��x	L	��h	L	��\	L	k�                	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~                         _., .   _   ;   C   =;  1#QNAN  1#INF   1#IND   1#SNAN  united-states   united-kingdom      trinidad & tobago       south-korea     south-africa    south korea     south africa    slovak  puerto-rico     pr-china    pr china    nz  new-zealand     hong-kong   holland     great britain   england     czech   china   britain     america     usa us  uk  swiss   swedish-finland     spanish-venezuela       spanish-uruguay     spanish-puerto rico     spanish-peru    spanish-paraguay    spanish-panama      spanish-nicaragua       spanish-modern      spanish-mexican     spanish-honduras    spanish-guatemala       spanish-el salvador     spanish-ecuador     spanish-dominican republic      spanish-costa rica      spanish-colombia    spanish-chile   spanish-bolivia     spanish-argentina       portuguese-brazilian        norwegian-nynorsk       norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg       german-lichtenstein     german-austrian     french-swiss    french-luxembourg       french-canadian     french-belgian      english-usa     english-us      english-uk      english-trinidad y tobago       english-south africa        english-nz      english-jamaica     english-ire     english-caribbean       english-can     english-belize      english-aus     english-american    dutch-belgian   chinese-traditional     chinese-singapore       chinese-simplified      chinese-hongkong    chinese     chi chh canadian    belgian     australian      american-english    american english    american        �	ENU �	ENU x	ENU h	ENA \	NLB P	ENC L	ZHH H	ZHI <	CHS (	ZHH 	CHS �	ZHI �	CHT �	NLB �	ENU �	ENA �	ENL �	ENC p	ENB `	ENI L	ENJ <	ENZ  	ENS  	ENT �	ENG �	ENU �	ENU �	FRB �	FRC �	FRL �	FRS l	DEA T	DEC <	DEL ,	DES 	ENI 	ITS  	NOR �	NOR �	NON �	PTB �	ESS �	ESB |	ESL h	ESO P	ESC 0	ESD 	ESF 	ESE �	ESG �	ESH �	ESM �	ESN �	ESI �	ESA p	ESZ `	ESR H	ESU 4	ESY 	ESV 	SVF  	DES �	ENG �	ENU �	ENU                                                                                                         �	USA �	GBR �	CHN �	CZE �	GBR �	GBR �	NLD �	HKG �	NZL �	NZL x	CHN l	CHN \	PRI T	SVK D	ZAF 4	KOR $	ZAF 	KOR �	TTO �	GBR �	GBR �	USA �	USA                                     6-    OCP ACP Norwegian-Nynorsk       C O N O U T $       ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               RSDSp�yoG}C�vC��?   C:\Program Files\MAXON\Cinema 4D R14.025\plugins\_Container Object\containerobject.pdb                                                                                                                                                                                                                                                                                                       @	|	               �	    �	�		T	     @	       ����    @   |	        $@	       ����    @   �	                    	    �		T	    D@	       ����    @   4	                   H	    	T	    `@	        ����    @   x	                   �	    T	                $@	�	                D@	4	                �@	�	               �	    �	    �@	        ����    @   �	                    �@	4 	               H 	    T 	�	    �@	       ����    @   4 	                    �@	� 	               � 	    � 	    �@	        ����    @   � 	                    A	� 	               � 	    !	�	    A	       ����    @   � 	                    $A	D!	               X!	    h!	!	�	    $A	       ����    @   D!	                    PA	�!	               �!	    �!	    PA	        ����    @   �!	                    `@	x	                �A	"	               ("	    0"	    �A	        ����    @   "	                    �A	l"	               �"	    �"	    �A	        ����    @   l"	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ����    ����    ����    ��    ����    ����    ��������    ����    ����    ����    ��    ����    ����    ����    `	    ����    ����    ����    k
    ����    ����    ����        ����    ����    ����    ~    ����    ����    ����        ����    ����    ����    �����    �        ����    ����    ����    �����    �        ����    ����    ����    �'    ����    ����    �����_�_    ����    ����    ����    �}    ����    ����    ����    ��    ����    ����    ����    Z�    ����    ����    ����    -�    ����    ����    ����    ��    ����    ����    ����    ג    ����    ����    ����    &�    ����    ����    ����    m�    ����    |���    ����    �    ����    |���    ����    F	    ����    ����    �����&�&    ����    ����    �����& '    ����    ����    ����    �'    ����    ����    ����    �*    ����    ����    ����    �,    ����    ����    �����/�/    ����    ����    ����    j=    ����    ����    ����    3G    ����    ����    ����    K    ����    ����    ����    �n    ����    ����    ����    �o    ����    ����    ����    �p    ����    ����    ����    2x����    >x        ����    ����    ����    y����    *y        ����    ����    ����    b�        �        1�            ����    ����    ����    7�    ����    ����    ����    ,�        h�        ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��        V�        ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    �2    ����    ����    ����    �3    ����    ����    ����    �l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���P    R0	          H0	 L0	 P0	 F� f0	   containerobject.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                  4�    .?AVContainerObject@@       4�    .?AVObjectData@@        4�    .?AVNodeData@@      4�    .?AVBaseData@@      8   �   �   �   �   �  �  c  �  4�    .?AVGeDialog@@      4�    .?AVGeModalDialog@@         4�    .?AVGeUserArea@@          �  4�    .?AVSubDialog@@     4�    .?AViCustomGui@@        w  �  �  4�    .?AVNeighbor@@      B  Q      (   2   4�    .?AVC4DThread@@     D   g   �   )      4�    .?AVtype_info@@     u�  s�              cos             asin            sqrt            N�@���D        ����������        ��������        �����
                                                                                                           	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                             ?     ��   ��   ��   ��   d�   \�!   T�   ��   ��   ��   L�   D�   ��   ��    ��   ��   ��   <�   ��   4�   ,�   $�   �   �"   �#   �$   �%    �&   ��                                                      �      ���������              �               �D        � 0                    ����                                                                                                                                                                                                                                                                                                                                        abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     �E	�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                            ����C   �����������������������������������������������t�l�d���\�T�L�@�4�(���������	         ����������������p�\�D�,�������������������������t�`�H�8�(����� �������������|�L�4�                                                                                                                                                                   L	            L	            L	            L	            L	                              8T	        �	@
	�	 L	                                            �M	�M	�E	        �p     ����    PST                                                             PDT                                                             �N	8O	                                ����        ����                                                                                                                                                                                                                                                                                                                                                                  �&       s	     s	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     .   .   0T	�o	�o	�o	�o	�o	�o	�o	�o	�o	4T	�o	�o	�o	�o	�o	�o	�o	8T	                    �	�	    ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                      �	     �                   ���5      @   �  �   ����                            .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                            ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (�	         ,�	 ̑	                     p�	 ��	 ��	 ��	 ��	 ̓	 ؓ	 �	 ��	 �	 �	 2�	 N�	 Z�	 h�	 v�	 ��	 ��	 ��	 ��	 Ԕ	 �	 ��	 �	 �	 "�	 2�	 Z�	 h�	 z�	 ��	 ��	 	 ؕ	 �	  �	 �	 (�	 8�	 N�	 Z�	 f�	 |�	 ��	 ��	 ��	 ޖ	 �	 �	 �	 �	 $�	 6�	 P�	 h�	 x�	 ��	 ��	 ��	 	 З	 �	 ��	 �	 �	 *�	 :�	 P�	 b�	 r�	 ��	 ��	 ��	 ��	 И	 ޘ	 �	  �	 �	                                                                                                         p�	 ��	 ��	 ��	 ��	 ̓	 ؓ	 �	 ��	 �	 �	 2�	 N�	 Z�	 h�	 v�	 ��	 ��	 ��	 ��	 Ԕ	 �	 ��	 �	 �	 "�	 2�	 Z�	 h�	 z�	 ��	 ��	 	 ؕ	 �	  �	 �	 (�	 8�	 N�	 Z�	 f�	 |�	 ��	 ��	 ��	 ޖ	 �	 �	 �	 �	 $�	 6�	 P�	 h�	 x�	 ��	 ��	 ��	 	 З	 �	 ��	 �	 �	 *�	 :�	 P�	 b�	 r�	 ��	 ��	 ��	 ��	 И	 ޘ	 �	  �	 �	                                                                                                          IsDebuggerPresent �GetCurrentThreadId  � DecodePointer �GetCommandLineA � EncodePointer �HeapAlloc GetLastError  �HeapFree  �GetTimeFormatA  �GetDateFormatA  yGetSystemTimeAsFileTime IsProcessorFeaturePresent �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �InterlockedIncrement  GetModuleHandleW  sSetLastError  �InterlockedDecrement  �GetCurrentThread  EGetProcAddress  �Sleep ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW WideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId �HeapSize  %WriteFile GetModuleFileNameW  �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter �RaiseException  GetLocaleInfoW  rGetCPInfo hGetACP  7GetOEMCP  
IsValidCodePage �GetTimeZoneInformation  9LeaveCriticalSection   FatalAppExitA � EnterCriticalSection  RtlUnwind �HeapReAlloc -SetConsoleCtrlHandler bFreeLibrary �InterlockedExchange ?LoadLibraryW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  -LCMapStringW  gMultiByteToWideChar iGetStringTypeW  �SetStdHandle  $WriteConsoleW �GetUserDefaultLCID  GetLocaleInfoA  EnumSystemLocalesA  IsValidLocale � CreateFileW R CloseHandle WFlushFileBuffers  d CompareStringW  VSetEnvironmentVariableA KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ,   �7�8�8\9�9�9":@:�:�:�:I;�;�;v<�<�<�? 0 H   22222 2$2(2,2�233�3�3�3436D6U6F9�9:B:�:�:	<�<�=�>�?�?�?   @ H   G0�081�1�1�1�1.2C23V3�3�3�3h4Q5f5�5_6q7�7
8�89/:f:"<b<�<=�>�? P �   �0�021r1�1�122v2�2�2"3]3�3�3�324~4�45f5�5�56b6�6�6.7v7�7�768y8�89i9�9":]:�:�:;E;z;�;�;9<z<�<�<I=�=�=>�>�>"?f?�?�?   ` @   >0}0�0�2�2�2�2�2�2�2�2333&303:3D3N3X3�4�7�<`>d>h>l>p> p    �0�0�0�<	=y= � L   �0F1�1�1	2N2�4�4F9}9�9_;n;};�;�;=<�<�<�<�<�<�<�<�<>_>�>�>#?Z?�?�?   � �   �0�0�0;1a1�1�1'2N2�2�2�2/3[3�3�34D4�4�455c5�5�5�56"66�6�67:7q7�7�7*8a8�8�8B9�9�9:U:�:�:2;~;�;<f<�<�<F=�=
>n>�>�>2?r?�?�? � 4   60y0�0;1�1�1�1�1�4�4�4�4�5�5
8A8�8�8"9i9�<   � H   �0�0�0�1�1�1�2�263�3�3
4:4j4�4�4V5�5�566y6�67R7�7�78U8�8%>�>�? � |   z0�0�0*1C1�1�12F2�2�23B3�3�3&4�425r5�5�566�6�67_7�7�768�8�8�8/9n9�9�95:m:�:�:&;h;�;�;<=<r<�<�<2=r=�=�=2>r>�>�>   � `   �3�3�3�4-626@67Y7�7#8c8�8�8&9b9�9�9$:Z:�:�:O;�;�;�;-<b<�<=I=�=�=�=>M>}>�>�>"?v?�?�?   � |   30v0�0�031s1�1�23O3�3�3&4_4�45E5R56�6�67F7z7�7�7=8m8�8�8"9b9�9�9":b:�:�:";b;�;�;"<b<�<�<"=b=�=�=&>f>�>�>I?�?�?   � t   0S0�0�01V1�1�12V2�2�23R3�3�34R4�4�45b5�5�5>6�6�6�627r7�7�7&8]8�8�8�8K9�9�9�<�<�<�<4=�=�=�>�>?X?�?�?     8   70{01v1�1	2r234c4�4D5�56z6�6:7�:�;�>�>�?�?�?  $   00�01�123�4f5�7�8:�<s=   H   0R0a0i162�2'3�34�45�56�67n7�7g8�8g9�9e:�:e;�;g<�<W=�=U>�>�? 0 \   U0�021�1�1J2�23E3�34�4�455S5�5	6v6�6>7�78�89�9�9a:�:�:8;�;�;G<�<�<W=�=>q>�>�?   @ l   �0�2�3�3�3�3�3�3�3�3�3�4�5 66666666�7a8w8�8!9@9`9�9�95:u:�:;t;�;=<B<�<�<=X=�=�=6>�>�>9?�?�? P \   0e0�182}2�23U3�3�3=4�45>5P5U5�5�5�5�566�67d7�7�748�8�8-9}9�92:�:?;�;�;<�=�>�? ` $   I2�2�3�3F4�4�5B66�9�9!:m:�: p     �0r1�1�1R2�23�3�3�;�?   � $   3�3�3�4�45=5u5�5�5�6�6�:   � d   2[2�2�23Y3�3�364t4�4�485t5�5�5I6�6�6�78V8�8�8)9y9�9:B:�:�:	;^;�;�;2<y<�<=N=�=�=>�>&?�? � l   G0�0
1?1�1�12r2�2�2f3�3�324r4�4�4b5�5�5;6�6�6"7z7�748q8�:�:�:�:�:;D;I;];�=�=�=�=	>>	?�?�?�?�?�?�? � 0   +303C3z33�3�4�4_5d5�6�6�6�6-:i:�:b?�?�? � P   0F0�0�0	1R1�1�12u2�2�2�3�3�34r4$5o5�56w6�67y9�9�;7<r<�<�>�>?Q?�?   � P   V0�01Q1�1�12V2�2�293�3�34^4�4�4&5f5�56}6�627v7�7�7�8�8 9969=7>�?   �    �1z5;y; �    �<a>�>}?�?�?   t   =0s0�0�0&1c1�1�12S2�2�223�3�3:4�4�445t5�5Y6�6�6r7�798�829r9�9
:A:z:�:�:I;�;�;<j<�<�<N=�=�=.>v>�>?C?�?�?�?  �   G0�0�01J1z1�1�1/2o2�23J3�3�3�3@4g4�4�45:5o5�5�56?6v6�6�6C7�7�7#8c8�8�8*9c9�9�9':z:�:�:c;�;�;6<v<�<�<6=s=�=�=/>o>�>?~?�?   \   :0�061�1�12r2�2�2!3_3�3�3
4?44�45_5�5�6�6&7�7�78_8�8�8^9�9:o:�:�:�:v;{;�;/<�?�? 0 |   0Y0�0�0&1f1�1�12g2�2�23_3�3�34f4�4�4&5_5�5�56Z6�6�6
7F7�7*8f8�89Y9�9�9>:�:�:&;Z;�;�;N<�<�<=^=�=�=N>�>?_?�?   @ �   0b0�031�1�2�2)3y3�3�455h5w55�5�5�5�5�566J6R6d6l6�6�6�6�6�6�6�6:7q7�7�7"8i8�8�8-9b9�9�9!:i:�:	;B;�;�;<V<�<�<2=r=�=>I>�>�>&?f?�?�? P 0   &0f0�0�021r1�1�192x2�2�2835�6B8:B:�:�: ` D   90�46�6�6*7a7�7�7!8�8�8W9�9�9:f:�:�:.;e<�<�=B>�>�>?F?�?�? p p   0O0T0Y0^0�0�1�1R2�2�23F3�3�34r466s6�6�67V7�7�7:8�8�8�8�89	9%9�9�9::�:�:I;N;;<K<o<<=�=!?0?9?>?D? � |   10G0�0�0A1z1�1�12�2�2l3�3�3�3�34)4�455�5�56B6�6�67v7�7\8�8�869v9�9�99:q:�:�:!;a;�;�;<T<�<�<=Q=�=�=�=�>?A?q? � X   "0b0�0�0"1b1�1�1"2b2�2�2"3b3�3�3"4b4�4/747E7o7t7�7�8�8�8�8�89):.:?:r:w:�:�:�:�: �    Z6   �    �7�7:   � x   �0<1@1D1H1L1�2�2"3b3�3�3&4b4�4�425v5�5�566r6�6�6�8�8�8�8O9p9�9�:�:;5;<<A<J<O<T<�<�<2>O>T>e>�>�>�>1?>?�?�?�?�?�? � �   !0A0q0�0�0�12v2�2	3#3^3I4�4�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�566R6n6(7`7e7o7�7�7�7�7898?8E8Z8�899l9�9J:Q:Y:�:�:�:�:6;;;@;c;�;r<�<='=9=D=q=|=�=�=2>�>�>�>??+?�?�?   �   "0-0?00�0�0�0111�1�1�1�1,2D2K2S2X2\2`2�2�2�2�2�2�2�2�2�2�2�2:3@3D3H3L3�3�3�3�3�3�3�3474i4p4t4x4|4�4�4�4�4�4�4�4�4�46Z6s6�677"7�7�7�7�7888898_8}8�8�8�8�8�8�8�8�8�8�8�8�8�8b9m9�9�9�9�9�9�9�9: :$:(:,:0:4:8:<:�:�:�:�:�:o<�<q={=�=�=�=�=�=�= >>\?d?y?�? �    �;N<U<>2>     (   *7�89!9�9�9�9�:�:�:V;[;�;�;�<    l   �071�1�8�9�;�;�;E<J<Y<b<u<{<�<�<�<�<�<�<�<�<�<�<=	===#=)=E=O=U=_=�=�=�=)>/>Y>_>e>{>�>�>W?z?�?�?�?      [0k0q0}0�0�0�0�0�0�0�0�0�0�0	1111#1)10161>1E1J1R1[1g1l1q1w1{1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122-232K2�2�2�2 3%3.3:3�3�3�3�3�3�3H4Q4]4�4�4�4�4�4�5�5�566%6*6<6F6K6g6q6�6�6�6�6�6�6�67D7N7t7{7�7�7�7�8�8�8(9m9t9�9�9�9::;:_:�:�:�:�:�:�;�;�;<<I<S<�<�<�<�<�<=4?E?M?S?X?^?�?�? 0 �   0B0�0�0�0�0�0131?1O1U1[1g1q1�1"2�23373�3�5!6.6:6B6J6V66�6�6�6�7�7 88I8U8e8q8�8�8�8�899�9Y:�:h;�;�<�=�=�=�=�=�=�>�>?d?q?�?�?�?   @ �   50F0�0�0�0�0�0�0I1U1]1�1�1�1#2R2Z2b2�2�3�3�3�5�5�526J6T6o6w6}6�6�6�6�67/7{78M8i8�8�8�9�9�9�9�9�9:::�;�;�;�;�;�;�;�;J<�<�<�<�<�<==:=C=L=b=�=�=�=�=�=�=�=�=�=�= >	>P>T>X>\>`>d>h>l>p>t>x>|>�>H?�?   P |   Q0W0]0c0i0o0v0}0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111"1(1>1E1�36636I6Q6�68*8�8�8I9�9C:�:?;�;�>�>�>9?Y?f?t?�?�?   ` H   0#0G0�01u1
22&282H2T2�34!4;4�4T5�5O6\7c7g9�9:C:�:�:�:>?   p t   V0�0�0�0�2�4�4�4�4�4�4�45�78�8�899�9�9�9�9�9�9�9::s:z:;Z;q;E=V=�=�=�=�=�=�=%>0>:>S>]>p>�>�>?2?�?�?   � �   0w0]1�1�1�122&2.2E2^2z2�2�2�2�2�2�2\3m3�3�3F4�45�5�5�6�67:78U8�8 9Y9_9e9k9�9":+:1:6:N:h:�:�:�:�:�:�:�:�:�:;;;(;H;R;�;�=�=�>�>�>�>�>?	???7???I?V?^?d?j?   � \   ,040@0M0T0\0d0l0u0~0�0�0�0�0�0�0�0�0�0�0�0X1]1�1�1I2V2i2v2�2�24::�=�=�?�?�?�?�?   � �   00<0C0\0�0�0�0�0�0�0.1�1�1E2e2�2�2�2�2�2'3f33�4�456C6S6_7}7�7�7�7�7�7�7�7�7�8�8�8	99+9<9R9c9t9�9�9�9�9�9�9�9�9>:P<c<�<E=v=~=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=)>@?F?W?]?f?m?t?}?�?�?�?�?   � `   0M0�0�1�12R2�2�3�3K4v4�4J5w5�647�739�9:-:�:;;�;�;3<�<�<�<=-=<=[=�=
>>?,?2?a?�?�? � �   �0�0�0�0�0�011)1w1{11�1�1�1�1�1�12+212=2D2h2z2�2�2�2�2�2�23,3U3�3�3�34y4�4�4�4�4;5B5M5�5'6@6Q79T9b9i9�9�9�9�9::�:�:�:�:�:�:�:;%;};�;�;�;�;�<�<�<= =�=�=�=�=>�?�?�?�?�?   � �   0C0�0�0111D1K1m1r1�1�1�1�12/2L2�2�2�2a3�3�3�3n4�4�4�475v5�5�5�5 66M6Z6�6�6�6�6�7>8]8m8z8�8�8�8�8�89�:�:�:�:�:�:;	;;N;�;�;�;�;�;U<a<{<�<�<�<�<�< ='=Q=c=�=�=�=�=>>4>"?6?a?m?�?   � l   0>0S0u0|0�0�0�0�011q1�1�1�1.2G2�3f4�4�4�4,6^6�6787P7�7K8�8�89G9:�:�:=;�;3<�<r=�=�==>�>�>�>?   � t   �2�2�2�2�2�2�283e3y3�3�3�3b4�4�4�5�5�5�5'676�6�6�6�6J7\7|7�7�78�829I9�9�9W:n:t:�:H;�;@<\<�=>P>�>�>a?f?�?�?   �   �0�0161N1[1�1�1�4�4585=5^5j5}5�5�5�5�5�5�5�5Q6�7�7�7'8/858;8A8h8�8�8�8�8�89(9{9�9�9�9�9�9�9�9�9/:7:s:�:�:�:�:�:�:;;;B;I;q;�;�;�;�;�;<<K<�<�<�<�<===!=%=)=1>p>�>�>�>�>�>?"?F?Y?�?�?�?�?�?  P   Y0�0�0�0�0�0U1�123:4F4�4�4y5�56#6�6�6\7h7�78�8�8E9Q9�9�9�:�:�<4=">?   �   00502�4�4�4T5Z5f5�5�5}6�6�6�67%7*7<7A7F7K7[7v7|7�7�7�7�7%8a8g8�8�8
9!9a9�9�9�9�9�9�9�9:	:::%:*:2:8:F:K:S:Y:g:l:X;�;�;�;�;�;�;�;�;	<j<s<y<i={=�=�=�=�=�=�=>#>+>9>X?]?o?�?�?�? 0 d   �3�485[5f5l5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�56<6V6p6;9B9H9{9�9�:�:E;(<5<N<�<�<�<�=>�>�>�?�?   @ d   R0�1�2j3�3�3�34m6�6�6z7�78:8@8Z8i8v8�8�8�8�8�8�8�8#919N9X9~9�9�9�9	:G:�:�;<<%<0<I=g=�?�? P    z0J1N2q2
3   ` `   2t2�233'393�3�4�4�4�4�4 5!636E6W6i6{6�6�6�6�6�6�6�6r7�9X:i:�;�;�;�;�;�;}<�<�<�<�>)?   p `   )0;12�3�4�4�4�4�5�5$6,6S6[6�6�6�6�647V7b7n7y7�7�7�78�89:�:H;j;�;�;�; <<<W<h<�<o=�=�> � H   02L2�2�2�2 4�4�4�4517�7�8�8�8�8�8�899�9:�:a;m;�;�;<a=m=   � ,   �0�7899�9�:B;H;�;�;�;�<�<>>�>�?�? � (   n0O1�1�1�2�2�2>3U3�4t6�9�9�9K=�= � 4   �0�0�3�3�3�3�344
44444�5�6�7�7�7�7D8h8 �    >2�6N:�< � h   �0�4�6�6747�7�7�7�7N8v8�8�8�89*99�9�9�9�9-:R:_:�:�:�:�:�;�;�;=<�<�<=*=K=9>�>?>?G?n?{?�?�?   � <   �0�0�01\1�1w2�2B3�34<4_4�4�4�7�7�7�7z;�;�;�;^=m=�? � D   
00;0d0x0�041p12u2�2�4�4�5�56!6|6�6�6"7l7u7�7�7�7"818�>     H   �=�=�=�=�=�=�=�=�=>>
>>>>>>">&>*>.>2>6>:>>>B>F>J>N>R>V>Z>     �7     H   D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 0 <   �1�1�1�1�1�23E3e3�3�325�5�56r6�6�6:�:9<|<�<�<�>   @ (   �0�0�0�0�0�0�0�0�67:7`78/8 9p? P ,   �1222S2V6�6D9H9L9P9T9X9\9`9M>?w?   ` <   �0�2�2/3?3,424>4M4�4�4�4�45A5f5�5�79;v;�;�;�;<B<   p �   0
0000"0(0.040:0@0F0L0R0X0^0d0j0p0v0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 111111$1*10161<1B1H1N1T1Z1`1f1l1r1x1~1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12o2�2 �    �2   � d   11111(4,4044484H7L8@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � ,  80<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4 555555 5$5(5,5054585<5@5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6074787�7�7T9X9\9`9d90;4;<;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;   � 4   T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � �   �1�1�=�=�=�=�=�= >>>>>>>> >$>(>,>0>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?�?�?�?�?�?�?�?�?�?�?�?�?�?  	 4    00000�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> 	 �   �5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7 8(80888@8H8P8X8`8h8p8x8�8�8�8�8�8�8�8�8�8�8�8p>t>�>�>�>�>�>�>�>�>�>�> ????(?@?H?L?T?l?�?�?�?�?�?�?�?�?�?�?�?    	 �   0(0,0@0H0L0T0l0�0�0�0�0�0�0�0�0�0�0 11 181<1P1X1\1`1h1�1�1�1�1�1�1�1�1�122 2(202H2`2d2x2�2�2�2�78808P8p8�8�8�8�8�8 9,9P9l9p9�9�9�9�9:0:P:p:�:�:�:�:�:�:;0;P;l;p;�;�;�;�;<0<P<\<�<�<�<�<�<�<==@=`=�=�=�=�=�=>0>P> @	 @   0$0D0`0�0�0�01$1P1�1�1 2$2(2,2024282<2@2D2t4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45555$5,545<5D5L5T5�5�5: <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=(>8>H>X>h>�>�>�>�>�>�>�>�>x?|?   P	 8   (10184<4@4D4H4L4P4T4X4\4h4l4p4t4x4|4�4�4�4�4�4(5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    