MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$       ��/���A���A���A������A���@�ݲA�	t����A�f����A�	t����A�	t���A�	t����A�cY���A�cY����A�cY����A�Rich��A�                        PE  L �n
R        � !    b      a�     0                         �         @                   �f O   Tc <                            � `                                  �: @            0 �                           .text   e                        `.rdata  /7   0  8                @  @.data   �   p     N             @  �.reloc  "   �  $   R             @  B                                                                                                                                                                                                                                                                                                                                                                        ��  �`r3ĉ�$�  ��$�  S��$�  U��$�  W��$�  �|$�l$�\$�D$����  ����  ��rV���   j ���   j��$l  Q���Ћ�rj ���   �����   j�D$,P�͉t$ �ҋ��~t3�3ۅ�~[���    ��4l  ;D4,uA��4d  ��t6�|4$ t/��r���   �@�Ћ�r�����   �L4$�R��;���   C;�|��\$���L$u��|$��$�   tn��r�ϋ��   �@8�Ћ���tV�l$ ��    ��r���   �ϋR,�ҋ�r�t$���   S��ϋ��ҋЅ�t��rU���   �ʋ@D�Ћ���u�^_]�   [��$�  3��� �Ę  ��t$��r�\$���   ��4h  �@S�t4,���4�����$�  _][3�3���� �Ę  ����V�t$W����   �|$����   S���NO  �ϋ��EO  ��t��tP���c ��u[_^á�rh� ���   �΋@�Ѕ�tx��rh� ���   �ϋ@�Ѕ�t]��rV�@@�@,�Ћ�rW�I@�؋I,�у�����t5��t1��rh�  �A�ˋ@T�ЋЅ�t��rR�Ah�  �@D����[_�   ^�_3�^�������������V�*  ���C  ��t��t�   ^�3�^á�rQ�@�@��Y�V���x%  �D$t	V�  ����^� ��j�hd�    P��HSUVW�`r3�P�D$\d�    �l$l��u3��1  �L$,�QK  �D$,Pj hbyek�D$p    踮  ��r���@j ���   haqpi�L$4�Ћ��L$@���&  ��r�D$d�A�L$�@Q�Ѓ��D$Pj�D$l�0> ���L$DPj j��(  ����r�L$�@Q�@���D$h�Ѓ����\  �   �   ��E�j P�D$HP��  ���D$��uj��= P�D�  ���   ���u�  �����  ��rhD� ���   �ϋR�҅�t3��r�ϋ��   �@(�Ѕ�u��r�ϋ��   �@L�Ћ߉\$�  hD� �b �؃��\$��uj�>= P踪  ���  ��r�ϋ��   �@x�Ћ�rP���   �ˋB|�С�rh  ���   �ϋ@�Ѕ�tK��r�ϋ��   �@(�Ѕ�u5PSW������r�����   j ��,  S����jj j SW�������T�D$l    �
��$    �I ��r�ϋ��   �@(�Ћ�r�����   �ϋRL��j �t$p��SW���  �|$l����u��L$�'�  ����tK3ۋ�r���   �ϋ@(�Ћ�r�����   �ϋRL��j SW���l�  Wj,����  �ߋ���u��\$�D$P��  ��rj �@@S�@�Ѓ���j j j S�K�  Sj,���q�  j S���g�  j ��  ���   �j�/�  ��3��L$@�D$d �%  �L$,�D$d�����H  �ƋL$\d�    Y_^][��T� ��̋V�t$V�P��u^� W����  h  �D$�G ������u_^� �t$��j-���  jj j W�t$�����j W�t$(�������r�L$,���   �� �@x�Ћ�rP���   �ϋB|�С�r�t$�@@�@�Ћ�rP�I@W�A�С�r�L$���   ����,  j W�С�r�t$���   �ϋ@@��Wj,���'�  ��r�L$���   �@L�ЍD$P�y j �B�  ���   _^� ����̋L$��t/��  �Ѕ�t$��rhD� ���   �ʋ@�Ѕ�t�   @� 3�� ����j�hid�    P��VW�`r3�P�D$$d�    h�0jnh�rj�H  �����|$�D$,    ��t���   ��0�3���r�L$�@Q�@�D$0�����С�rj �@j��@�L$ h�0Q�Ѓ��D$P�L$�D$0   �P  �0Wj�D$4�E9 ��PVh   j�49 ��Ph:� �62 ���L$���D$,�R  ��r�D$�IP�I�D$0�����у��ƋL$$d�    Y_^��$��j�h�d�    P��VW�`r3�P�D$$d�    h�0h�   h�rj�%  �����|$�D$,    ��t����  �1�3���r�L$�@Q�@�D$0�����С�rj �@j��@�L$ h<1Q�Ѓ��D$P�L$�D$0   �qO  �0Wj
�D$4�"8 ��PVh   j	�8 ��Ph;� �1 ���L$���D$,��P  ��r�D$�IP�I�D$0�����у��ƋL$$d�    Y_^��$����������������K  �v����   ������������������L$t�   ù|r�Z5 ����������VW�|$3���t{S�\$$U�l$$��t
Wj0�����  �t$���t$�=G  ��r�ϋ��   �@4�ЋL$ ��t��tSUQ�t$(�t$(P��������t���r�ϋ��   F�R(�ҋ���u�][_��^�����VW�|$3���tGS�\$U�l$���$    ��t$���F  ;�uF��u��r�ϋ��   �@(�Ћ���u�][_��^�_��^���������V�t$j j�t$j?�t$������t$(��j j�t$0jP�t$4�������0��^���������j�h�d�    P��SUVW�`r3�P�D$(d�    �D$    ��r�\$8�@S�@�D$4    �С�r�l$@�@S�@U�Ѓ���r3��@�͋@<�D$0    �D$   �|$�Ѕ��0  �d$ ��rW�@S�@4�Ћσ��Ё�  �yI�ɀA��p����ȋ��ȉD$ ���(������D$$;���   �|$ ��$    ��r�L$<�@�@<�Ћȋƙ����r�@�@4R�t$<�Ћ΃��Ё�  �yI�ɀA��p��L$<D$��r�@�@<�Ћȋř���L$I��ك��;t$$|��|$��r�H��  �yK�ˀC��
f�Ë\$8��P�A8WS�Ћ�rG�Q�L$H�R<���|$��;�������ËL$(d�    Y_^][�� ���������������j�h,d�    P��$V�`r3�P�D$,d�    ��r�L$�@Q�@�С�rj �@j��@�L$(hX1Q�С�r�L$ �@Q�@�D$L    �С�rj �@j��@�L$,hh1Q�Ѓ�(�D$P�L$�D$8�K  h�  �0�D$Ph� j j �D$L�3 ��PhD� ��� ���L$���D$4�L  ��r�D$�IP�I�D$8 �ѡ�r�L$ �@Q�@�D$<�����Ѓ��ƋL$,d�    Y^��0�������������V���HE �F    �F    ��^������̡�rV���   �񋀌   V�Ѓ��    ^��������������̋	���f�  �������G ������������;  �����������j�hXd�    PQV�`r3�P�D$d�    ��t$��r�D$    �P�FP�B�Ѓ����D$������  �D$t	V�   ���ƋL$d�    Y^��� ��������j�h�d�    PQV�`r3�P�D$d�    h�2h�   h�rj �x  �����t$�D$    ��t:���L  �2��r�D$�Q�NQ�J�у��ƋL$d�    Y^���3��L$d�    Y^���������SUW�t$ �|$�t$ ���t$ �t$ W��F  ���u_][� � V�wt	V�u_ ���K��t��Z ��C�G��r�H�GP�CP�A�Ѓ���^_][� �������������V�t$���4F  ���> t	V�_ ��^� ���������������j�h�d�    P��SVW�`r3�P�D$ d�    ���|$0 �  �t$4���  hD� ���L ����   ��r���   ���   �ЉD$0h�  �L$�D$,    �C �t$0�D$P���D$0�[M �L$���D$( ��D h�  �L$��B �t$0�D$P���D$0�(M �L$���D$( ��D ��t��r�w�Aj�@0���Ѕ�t��r�w�@j�@0���ЋD$8�L$0���rQ���   �D$,�������   �Ѓ��   �L$ d�    Y_^[��� 3��L$ d�    Y_^[��� ������������j�hd�    P��(SVW�`r3�P�D$8d�    ���t$HV�^D  �؅�u�L$8d�    Y_^[��4� ��rV�@@�@,�Ћ�r���Q���R4jh�  ������2��r�D$ ��2�D$(��2�D$0�@�L$ �@HQh�  ���Ѓ �Gt	P��\ ���G    ��r�L$�@Q�@�С�rj �@j��@�L$h�2Q�С�r�O�@Q�@�L$(Q�D$\    �С�r�L$,�@Q�@�D$`�����Ѓ� �ËL$8d�    Y_^[��4� ��������������j�h�d�    P��VW�`r3�P�D$ d�    �t$4�D$    ��r�L$�@Q�@(�Ћ���r�|$8�IW�I�D$4   �ѡ�rW�@V�@�Ћ�r�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� �����������S�\$U�l$V�t$WUVS���B  �D$��u_^][� ��Ft1��t��uKS���~  �D$_^][� US���:   �D$_^][� S����
  �D$_^][� ���F u	US���{  �D$_^][� j�hXd�    P��HSUVW�`r3�P�D$\d�    �١�r�t$l���   �΋@T�Ћ��|$l��t�����  �L$pj �D$h    ��A � /������g  �$�D( �{ �V  Wj���R�  P�����ؽ�  �n�{ �3  Wj��3��-�  P������  �K��r�΋��   �@4��WjP�u������'�{ ��  ��rW���   j�@4��3���P�J�����  ����t
Vj*���d�  ��rV�@@�@,�Ћ��D$SP������P��rU�A�΋@8�D$l�С�r�L$�@Q�@�D$h ���j  �{ �c  �L$$�  �D$@jP�D$l�6  ��P�L$(�D$h�  �L$@�D$d�O  ��r�L$�@Q�@�Ѓ��D$Pj�D$l��* ���L$(Pj j�  ��r���I�D$�IP�D$h�у�����   �K����u	��X ���T ���u#j�* P��  ���L$$�D$d �  �   j j��D$,P�$U ��t j���  S�X ���L$$�D$d �  �Y�ZX j j��j@j@���	U �jjh   V�hU S�BX ���3�L$$�D$d �?  ��{ u���; t	S�X ���D$d������t���s�  �L$\d�    Y_^][��T� � & & ( �% �% ( ( �& ( ��������j�h�d�    P��\SVW�`r3�P�D$ld�    �ٍL$X�6  �D$XPjhbyekǄ$�       胙  ������  ��rj �@haqpi���   �L$`�Ш��  ��r�|$|���   �ϋ@T�Ћ���t���r�  Wj*����  ����  �{ ��r�@�@��  �L$(Q�ЍD$,P�D$|�V�  ����tl��r�L$8�@Q�@�ЍD$<P�D$|�.�  ����t*��r�L$8�@Q�@x�L$,�Ѕ�tFj�v( P��  ����r�L$8�@Q�@�D$x�Ѓ���r�L$(�@Q�@�D$x ���  �L$�����h�  �L$�D$x��: �D$P�L$�D$x��= �L$�D$t�< ��r�L$���   Q�@j����h�  �L$�: �D$P�L$�D$x�= �L$�D$t�r< ��r�L$���   Q�@j���ЍD$(P�D$LP�J����C   ��r�K�@Q�@�L$TQƄ$�   �С�r�L$X�@Q�@Ƅ$�   �Ѓ��L$�D$t��; ��r�L$8�@Q�@�D$x�ЍL$,�X  �L$8Q�ЍD$<P�D$|��  ����u�D$t��r�L$8�@Q�@���S  �D$8P�D$LP��������r�T$H�@�K�@xR�D$x�Ѕ�tj�& P�%�  ����C    �L$�8 �D$     �D$$    h�  �L$�D$x	�9 �D$P�L$�D$x
�< �L$�D$t	�; ��r�L$���   Q�@j����h�  �L$��8 �D$P�L$�D$x��; �L$�D$t	��: ��r�L$���   Q�@j���ЍL$�D$t�: ��r�L$H�@Q�@�D$x�ЍL$<��rQ�@�D$| �@�С�r�����   j �@j����j ��  ���L$X�D$t�����2  �L$ld�    Y_^[��h� �����̃�X�ISUVW�|$p��\$4�3��tL��tV�O ���N ����rV�I�D$     �I�D$$    �ы�rV�I��I�D$�у��L��u�S j j��j@j@���O ShD� �~ ����t�V�N �C�k�D$�C�D$ �C�l$�D$����  ��r�t$l�@@�@,�Ћ�r���Q�����   j h�  ���҉D$$���  ��rW��L$8Q�D$<�D$D�D$L�@h�  ���   �L$XQ�����~ ��2�~P�~X�Y��Y��Y��,��ΉD$0�,D$,�,ÉD$(�P ��r�؋ř����   �L$l�R4���D$$�D$�ҋ�����   j?���3  ��t��r�ϋ��   �@(�Ћ���u��x   3�9l$~p�D$�L$��|^�|$ O|$�D$$�t$(��r�t$0�@�t$8��  WUV�Ѓ���t��rh�   �@W��  USV�Ѓ�O�L$$u��D$�L$E;�|��L$l��  ������   �d$ j?����2  ��t��r�ϋ��   �@(�Ћ���u��}   3�9l$~u�D$�L$��I ��|^�|$O|$�D$l�t$(��r�t$0�@�t$8��  UWV�Ѓ���t��rh�   �@U��  WSV�Ѓ�O�L$lu��D$�L$E;�|��\$4�D$�C�D$ �C�D$�C�D$_�3�C�D$l^]�@   [��X� �G    _^][��X� j�hd�    P�� VW�`r3�P�D$,d�    ��r�t$<�@@V�@,�Ѓ���j j jj?�����  P�����P�D$$P������P��rh�  �A�ϋ@8�D$<    �С�r�L$�@Q�@�D$8�����С�r�����   �΋@4��j j jj?P�v���P�D$4P�;�����P��rh�  �A�ϋ@8�D$<   �С�r�L$�@Q�@�D$8�����Ѓ��L$,d�    Y_^��,� ���������S�\$UVW�|$SW�t$���6  ���t;�D$P����#  ��t+�|$ t-�N��t�J ��N �F�v���Z$  ��u_^]3�[� �~ �Ft	P�N �����  |#�^S���#  ��t΃; t�FP����#  ��t�_^��][� �������SVW�|$W�t$���}5  ��3���t[9F����P�W!  ��u_^3�[� �F��tjj h�� P����!  ��t��v���%!  ��t΃~ t�FP���!  ��t���_^[� ���̋�r�D$��t�I�   ;�j B�j P���   �Ѓ�ù   ;�VB�W�xW��0������u_^�Wj V�� �������_�F�xr   ^ËL$��t,�=xr t�y���A�u
�D$�%�0��r�L$�@� �������������̋L$��t,�=xr t�y���A�u
�D$�%�0��r�L$�@� �������������̋�r�D$��t�I�   ;�j B�j P���   �Ѓ�ù   ;�VB�W�xW��0������u_^�Wj V�!� �������_�F�xr   ^Ë�r�D$��t�I�   ;�j B�j P���   �Ѓ�ù   ;�VB�W�xW��0������u_^�Wj V�� �������_�F�xr   ^Ë�r�D$��t�I�   ;�j B�j P���   �Ѓ�ù   ;�VB�W�xW��0������u_^�Wj V�A� �������_�F�xr   ^á�r�t$�@� ��Y��������������̡�r�t$�@� ��Y��������������̋L$��t��r�L$�@��@  �����̡�rhﾭދ@��@  ��Y����������V�t$���t��rQ�@� �Ѓ��    ^�������������̡�r�@���  ���D$��t�x��u�   �3����������̡�r�@��  �࡜r�@��   ����r�D$��t"�t$�I�t$�   ;�B�P���   �Ѓ�ù   ;�VB�W�xW��0������u_^�Wj V��� �������_�F�xr   ^������������̋L$��r�ɺ   Dʅ�t�t$�@�t$���   Q�Ѓ�Ã�VB�W�yW��0������u_^�Wj V�R� �������_�F�xr   ^�̡�r�t$�@� ��Y��������������̡�r�t$�@� ��Y��������������̋D$�   ;�VB�W�xW��0������u_^Ã|$ tWj V��� ��_������F�xr   ^�̋�r�D$��t<�|$ �t$�I�t$�   t;�B�P���   �Ѓ�Ã�B�P���  �Ѓ�ù   ;�VB�W�xW��0������u_^Ã|$ tWj V�,� ��_������F�xr   ^�����������̋L$��r�ɺ   Dʅ�t+�|$ �t$�@�t$Qt���   �Ѓ�Ë��  �Ѓ�Ã�VB�W�yW��0������u_^�Wj V�� �������_�F�xr   ^��������������̡�r�t$�@� ��Y��������������̡�r�t$�@� ��Y�����������������2������������2���������̅�t�j������̡�r�@��  �࡜r�@��(  ��j�hMd�    P�� �`r3�P�D$$d�    �D$    ��r�T$�@R��   �ЋL$4P�D$0   �  �L$�D$   �D$, �  �D$4�L$$d�    Y��,� �̡�r�@��$  �࡜r�@��  �࡜r�@���  �࡜r�@��  �࡜r�@���  �࡜r�@��x  �࡜r�@��|  �࡜r�@��d  �࡜r�@��p  �࡜r�@��t  ���D$V����2t	V��������^� ̡�r�@$�@X����̡�r�@$�@\������t$��r�t$�@$�t$�@`Q�Ѓ�� j�hxd�    PQV�`r3�P�D$d�    ��t$��rV�@�@�С�rV�@$�D$    �@D�Ѓ��ƋL$d�    Y^�����������������j�h�d�    PQV�`r3�P�D$d�    ��t$��rV�@�@�С�rV�@$�D$    �@D�С�r�t$$�@$V�@d�Ѓ��ƋL$d�    Y^��� ����������j�h�d�    PQV�`r3�P�D$d�    ��t$��rV�@�@�С�rV�@$�D$    �@D�С�r�t$$�@$V�@�Ѓ��ƋL$d�    Y^��� ����������j�h�d�    PQV�`r3�P�D$d�    ��t$��rV�@�@�С�rV�@$�D$    �@D�С�rV�@$�t$(�@L�Ѓ��ƋL$d�    Y^��� ����������j�hd�    PQV�`r3�P�D$d�    ��t$��rV�@$�D$    �@H�С�rV�@�D$�����@�Ѓ��L$d�    Y^����������̡�r�t$�@$Q�@L�Ѓ�� �������̡�r�@$�@����̡�rQ�@$�@�Ѓ����������������j�h@d�    P��VW�`r3�P�D$ d�    �D$    ��rQ�@$�L$�@Q�Ћ���r�|$8�IW�I�D$4   �ѡ�rW�@V�@�Ћ�r�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� � ����������̡�r�t$�@$Q�@�Ѓ�� ��������j�h�d�    P�� VW�`r3�P�D$,d�    �D$    ��rQ�@$�L$�@ Q�Ћ���r�|$D�IW�I�D$@   �ѡ�rW�@$�D$D�@D�С�rW�@$V�@L���D$$   ��r�L$(�@$Q�@H�D$P   �Ћ�r�D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,� ��������������j�h�d�    P�� VW�`r3�P�D$,d�    �D$    ��rQ�@$�L$�@$Q�Ћ���r�|$D�IW�I�D$@   �ѡ�rW�@$�D$D�@D�С�rW�@$V�@L���D$$   ��r�L$(�@$Q�@H�D$P   �Ћ�r�D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,� ��������������j�hd�    P�� �`r3�P�D$$d�    �D$P�D$    ������t$4���D$0   �(����D$   ��r�L$�@$Q�@H�D$0   �Ћ�r�D$�IP�I�D$4 �ыD$<���L$$d�    Y��,� ����̡�rQ�@$�@(��Yá�rQ�@$�@h��Yá�r�t$�@$Q�@,�Ѓ�� �������̡�r�t$�@$Q�@0�Ѓ�� �������̡�r�t$�@$Q�@4�Ѓ�� �������̡�r�t$�@$Q�@8�Ѓ�� �������̡�r�t$�@$�t$�@PQ�Ѓ�� ���̡�r�t$�@$Q�@T�Ѓ�� �������̡�r�@$�@l����̡�r�@$�@p����̡�rV�@$��@LV�t$�Ѓ���^� ��j�hXd�    PQV�`r3�P�D$d�    �D$    ��r�t$�@V�@�D$    �С�rV�@$�D$   �@D�С�rV�@$�t$,�@L�Ћ�r�t$4�I$V�I@�D$,    �D$    �у��ƋL$d�    Y^�������������̡�rV�@$�t$�@@��V�Ѓ���^� �̡�r�t$�@$Q�@<�Ѓ�� �������̡�r�t$�@$Q�@<�Ѓ����@� ��̡�r�@(�@����̡�r�@(�@����̡�r�@(�@����̡�r�@(�@����̡�r�@(�@ ����̡�rj�t$�@(�t$�@��� �������t$��r�t$�@(�t$�@$��� ���̡�r�@(�@(����̡�r�@(�@,����̡�r�@(�@0����̡�r�@(�@4����̡�r�@(�@X����̡�r�@(�@\����̡�r�@(�@`����̡�r�@(�@d����̡�r�@(�@h����̡�r�@(�@l����̡�r�@(�@p����̡�r�@(�@t����̡�r�@(�@x����̡�r�@(���   ��j�h{d�    P��V�`r3�P�D$d�    ��r�L$�@Q�@�Ѓ��D$P���D$$    �   ��u3����r�L$�@$Q�t$,�@�Ѓ��   ��r�D$�IP�I�D$$�����у��ƋL$d�    Y^��� ��������Q��r�T$�@(R�@X�Ѕ�uY� �D$3�8L$����   Y� �������������j�h�d�    P��V�`r3�P�D$ d�    ��r�D$    �D$    �@(�L$�@hQ���Ѕ���   �L$��r��uM�@�L$�@Q�С�r�t$4�@�L$�@Q�D$4    �С�r�L$�@Q�@�D$8�����Ѓ��   �@h�2���   he  Q�Ћȡ�r���L$�@(��u�@4j�����3��L$ d�    Y^��$� �@j �t$Q���Ѕ�u"�D$P�?�����3��L$ d�    Y^��$� ��rj �H�D$HP�t$�A�t$<�ЍD$P� ������   �L$ d�    Y^��$� ����̡�rV�@(W�|$�@pW���Ѕ�t8��r�΋P(�GP�Bp�Ѕ�t!��r�΋P(�GP�Bp�Ѕ�t
_�   ^� _3�^� ������̡�rV�@(W�|$�@tW���Ѕ�t8��r�΋P(�GP�Bt�Ѕ�t!��r�΋P(�GP�Bt�Ѕ�t
_�   ^� _3�^� ������̡�rS�@(V�@pW�|$W���Ѕ���   ��r�΋P(�GP�Bp�Ѕ���   ��r�΋P(�GP�Bp�Ѕ�tn��r�_�@(S�@p���Ѕ�tW��r�΋P(�CP�Bp�Ѕ�t@��r�΋P(�CP�Bp�Ѕ�t)�GP��������t�G$P��������t_^�   [� _^3�[� ��������̡�rS�@(V�@tW�|$W���Ѕ���   ��r�΋P(�GP�Bt�Ѕ���   ��r�΋P(�GP�Bt�Ѕ�tn��r�_�@(S�@t���Ѕ�tW��r�΋P(�CP�Bt�Ѕ�t@��r�΋P(�CP�Bt�Ѕ�t)�G0P���/�����t�GHP��� �����t_^�   [� _^3�[� ��������̡�r�@(�@8����̡�r�@(�@<����̡�r�@(�@@����̡�r�@(�@D����̡�r�@(�@H����̡�r�@(�@L����̡�r�D$�@(Q�@P�$��� ���̡�r�D$�@(���@T�$��� �̡�r�t$�@(�t$�@|��� ��������j�h�d�    P��V�`r3�P�D$d�    ��L$(�D$P�|���P���D$$    �\   ��r���I�D$�IP�D$$�����у��ƋL$d�    Y^��� ������̡�r�|$ �P(�����D$�B8������Q��rV�@W�@d���L$j �Ћ�rh�2�I�p���   h�  V�ыȡ�r���L$��u�@(j��@4����_3�^Y� �@j �@hVQ�L$�С�rV�@(�ϋ@H�Ѕ�t2��rV�@(�t$�@ ���Ѕ�t�D$P�   �x�������_^Y� �D$P3��a�������_^Y� �����̡�rV�@(W�|$�@P�Q���$�Ѕ�tF��r�G�@(Q�@P���$�Ѕ�t(��r�G�@(Q�@P���$�Ѕ�t
_�   ^� _3�^� ��rV�@(W�|$�@T������$�Ѕ�tJ��r�G�@(���@T���$�Ѕ�t*��r�G�@(���@T���$�Ѕ�t
_�   ^� _3�^� ���������̡�rV�@(W�|$�@P�Q���$�Ѕ��  ��r�G�@(Q�@P���$�Ѕ���   ��r�G�@(Q�@P���$�Ѕ���   ��r�G�@(Q�@P���$�Ѕ���   ��r�G�@(Q�@P���$�Ѕ���   ��r�G�@(Q�@P���$�Ѕ�ts��r�G�@(Q�@P���$�Ѕ�tU��r�G�@(Q�@P���$�Ѕ�t7��r�G �@(Q�@P���$�Ѕ�t�G$P���������t
_�   ^� _3�^� ��������̡�rV�@(W�|$�@T������$�Ѕ���   ��r�G�@(���@T���$�Ѕ���   ��r�G�@(���@T���$�Ѕ���   ��r�G�@(���@T���$�Ѕ�th��r�G �@(���@T���$�Ѕ�tH��r�G(�@(���@T���$�Ѕ�t(�G0P���T�����t�GHP���E�����t
_�   ^� _3�^� ��r�@(� �����̡�rV�@(�t$�@�6�Ѓ��    ^�̡�r�@(���   �࡜r�@(�@����̡�r�@(�@����̡�rV�@(�t$�@�6�Ѓ��    ^�̡�r�t$�@,�t$�@Q�Ѓ�� ���̡�r�@,�@����̡�r�@,�@����̡�r�@,�@����̡�r�@,�@ ����̡�r�@,�@(����̡�r�@,�@$����̡�r�@,�@�����j�hd�    P�� VW�`r3�P�D$,d�    �D$    ��r�T$�@,R�@�Ћ���r�|$<�IW�I�D$8   �ѡ�rW�@$�D$<�@D�С�rW�@$V�@L���D$   ��r�L$ �@$Q�@H�D$H   �Ћ�r�D$$�IP�I�D$L �у��ǋL$,d�    Y_^��,� ��������������̡�rj �@,j � �Ѓ�������������̡�rV�@,�t$�@�6�Ѓ��    ^�̡�r�@,�@4����̡�r�@,�@8�����j�hYd�    P�� VW�`r3�P�D$,d�    �D$    ��r�T$�@,R�@<�Ћ���r�|$<�IW�I�D$8   �ѡ�rW�@$�D$<�@D�С�rW�@$V�@L���D$   ��r�L$ �@$Q�@H�D$H   �Ћ�r�D$$�IP�I�D$L �у��ǋL$,d�    Y_^��,� ���������������j�h�d�    P��VW�`r3�P�D$ d�    �t$4�D$    ��r�T$�@,R�@@�Ћ���r�|$0�IW�I�D$,   �ѡ�rW�@V�@�Ћ�r�D$�IP�I�D$   �D$8 �у��ǋL$ d�    Y_^�� � �������̡�r�@,�@,����̡�rV�@,�t$�@0�6�Ѓ��    ^�̡�r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@�@����̡�r�@�@����̡�r�@�@����̡�r�@�@����̡�r�@�@����̡�r�@�@����̡�r�t$�@�t$�@\��� �������̡�r�t$�@�t$��  ��� ����̡�r�D$�@���@ �$��� �̡�r�D$�@Q�@$�$��� ���̡�r�D$�@���@(�$��� �̡�r�@�@,����̡�r�@�@0����̡�r�@�@4����̡�r�@�@8����̡�r�@�@<����̡�r�@�@@����̡�r�@�@D����̡�r�@�@H����̡�r�@�@L����̡�r�@�@P����̡�r�@���   �࡜r�t$�@Q��  �Ѓ�� ����̡�r�@�@T����̡�r�@�@X����̋T$��u3�� ��rR�@ Q�@(�Ѓ��   � ��������̡�r�@���   �࡜r�@�@`����̡�r�@�@d����̡�r�@�@h����̡�r�@�@l����̡�r�@�@p����̡�r�@�@t����̡�r�@���   �࡜r�@��  �࡜r�@�@x����̡�r�@�@|����̡�r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�t$�@Q��  �Ѓ�� ����̡�r�@���   �࡜r�@���   ���T$��t��rR�@ Q�@$�Ѓ���t�   � 3�� ����̡�rQ�@ �t$�@L�t$�Ѓ�� ���̡�r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜rV�@�t$���   V�Ѓ��    ^���������������̡�r�@� �����̡�r�@�@����̡�r�@���   �࡜r�@��   �࡜r�@�@����̡�r�@�@����̡�r�@�@����̡�r�@�@����̡�r�@�@����̡�r�@���  �࡜r�@�@�����j�h�d�    P��V�`r3�P�D$$d�    �t$4�D$P���|�����r�L$�@$Q�@�D$0    �Ѓ���t_��r�L$�@j�@Q�Ѓ���u�D$P��������t3��rj�@V�@�Ѓ���u��rV�@�@�Ѓ���t�   �3���r�L$�@$Q�@H�D$0   �Ћ�r�D$�IP�I�D$4�����у��ƋL$$d�    Y^��(���������������̡�r�@�@ ����̡�r�@�@(����̡�r�@��  �࡜r�@��   �࡜r�@��  �࡜r�@��  ��j�hd�    P�� VW�`r3�P�D$,d�    �D$    ��r�L$�@Q�@$�Ћ���r�|$@�IW�I�D$<   �ѡ�rW�@$�D$@�@D�С�rW�@$V�@L���D$    ��r�L$$�@$Q�@H�D$L   �Ћ�r�D$(�IP�I�D$P �у��ǋL$,d�    Y_^��,��j�hXd�    P�� VW�`r3�P�D$,d�    �D$    ��r�L$�@Q���  �Ћ���r�|$@�IW�I�D$<   �ѡ�rW�@$�D$@�@D�С�rW�@$V�@L���D$    ��r�L$$�@$Q�@H�D$L   �Ћ�r�D$(�IP�I�D$P �у��ǋL$,d�    Y_^��,���������������Qj�t$�D$    �  �D$�������j�h�d�    P��<SVW�`r3�P�D$Ld�    �D$    ��r��t�D$0P�.������D$T   �   �@��r�L$�@Q�@�С�r�L$�@$Q�@D�D$\   �Ѓ��|$�D$T   �   ��r�t$\�@V�@�\$�С�rV�@$�D$\   �@D�С�rV�@$W�@L�Ѓ�����t;����\$��r�L$�@$Q�@H�D$X   �С�r�L$�@Q�@�D$\�Ѓ��D$T    ��t<����\$��r�L$0�@$Q�@H�D$X   �Ћ�r�D$4�IP�I�D$\ �у��ƋL$Ld�    Y_^[��H���������������j�h*	d�    P�� VW�`r3�P�D$,d�    �t$@�D$    ��r�L$�@Q���  �Ћ���r�|$D�IW�I�D$@   �ѡ�rW�@$�D$D�@D�С�rW�@$V�@L���D$$   ��r�L$(�@$Q�@H�D$P   �Ћ�r�D$,�IP�I�D$T �у� �ǋL$,d�    Y_^��,����������̡�r�@��D  �࡜r�@��H  �࡜r�@��L  ��j�hf	d�    P��VW�`r3�P�D$ d�    �t$8�D$    ��r�t$8�@�L$���  Q�Ћ���r�|$<�IW�I�D$8   �ѡ�rW�@V�@�Ћ�r�D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� ���̡�r�@���  �࡜r�@���  �࡜rV�@j �@j����Ћ�^��������̡�rV�@j �t$�@���Ћ�^� ���̡�rV�@�t$�@j����Ћ�^� ���̡�r�@�@����̡�rV�@j ���   ��L$j V�Ћ�^� �������������̡�r�t$�@Q�@�Ѓ�� �������̡�r�t$�@Q�@�Ѓ����@� ��̡�rh#  �t$�@�t$�@l��� ��̡�rhF  �t$�@�t$�@l��� ��̡�r�t$�@�@t�Ћ�rP���   �@X�Ѓ�� ������̡�r�t$�@�@t�Ћ�r�t$�Ћ��   R�@`�Ѓ�� ̡�r�t$�@���   �Ћȅ�u� ��rQ���   �@�Ѓ�� �����������̡�r�@���   ���A    �    �A    �A   ������t$��r�t$�@@�t$�@Q�Ѓ�� ��r�t$�@@Q�@�Ѓ�� �������̡�r�t$�@@�t$�@Q�Ѓ�� ���̡�r�t$�@@Q�@ �Ѓ�� �������̡�r���   �@�࡜r���   �@�࡜r���   �@ �࡜r���   �@$�࡜r���   ���   ��������������̡�r���   ��D  ��������������̡�r�t$�@@Q�@L�Ѓ�� �������̡�rQ�@@�@H�Ѓ���������������̡�r���   ���   ��������������̡�r���   ���   ��������������̡�rQ�@H���   �Ѓ�������������V��L$��t2�T$��r���   ��t
�@@R��^� �T$�@D��tR��^� V��^� ��������������̡�r�@@�@0�����V�t$���t��rQ�@@�@�Ѓ��    ^������������̡�rV�@@��@V�ЋЋD$����t��#��С�rR�@@V�@�Ѓ�^� �����t$�D$��r�����   �$�t$���   �t$�t$�t$��� �������̡�r���   ���   ��������������̡�rQ�@H���   �Ѓ������������̡�r�t$�@HQ��d  �Ѓ�� ����̡�r�@@�@T����̡�r�@@�@X����̡�r�@@�@\����̡�r�@@�@`����̡�r�@@�@d����̡�r�@@�@h����̡�r�@@�@l����̡�r�@@�@p����̡�r�@@�@t����̡�r�@@�@x����̡�r�@@�@|����̡�r�@@���   �࡜r�@@���   �࡜r�@@���   �࡜r���   �@t�࡜r�@@���   �࡜r�@@���   �࡜r�@@���   �࡜r�@@���   �࡜r�@@���   �࡜r�@@���   �࡜r�@@���   ��V�t$���t��rQ�@@�@�Ѓ��    ^������������̡�r�@@�@0����̡�rj�@@�L$�@4Qj �Ѓ�������̡�rj�@@�L$�@4Qh   @�Ѓ����̡�r�t$�@@�t$�@4j �Ѓ������̡�r�@|� ������V�t$���t��rQ�@|�@�Ѓ��    ^������������̡�r�@|�@ �����V�t$���t��rQ�@|�@(�Ѓ��    ^������������̡�r�@ �@H����́|$qF uKW�|$��tA��r�t$���   �ϋ@D�С�r�t$�@@�@,�Ћ�r���ЋAW�t$�@p����_����������̡�r�@��T  �࡜rS�@@V�@,W�t$�Ћ�r�t$�I@�؋I,�ы�r���yh��hE  �ˋ��	���Ph��hE  �������P��T  �Ѓ�_^[�������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������3�� �����������3�� ����������̋L$�D$�A4�D$�A �D$��D$�A0�D$�A�8 �A8k �A<dO�A@sO�ADiO�AHnO�ALk �AP'k �Al,k �AX6k �A\;k �A`Ek �Ad@k �AT"k �Ah1k �ApJk �AtOk �A(�A,    �����������́�   h�   �D$j P��� j ��$�   �D$��$�   ��$�   ��$�   P������$�   h�   �D$T�D$(P��$�   ��$�   j�7�  ���   �j�h�	d�    P��   SV�`r3�P��$�   d�    ��� ����H  ��$�   �L$ ������r�L$�@Q�@Ǆ$�       �С�rj �@j��@�L$h3Q�Ѓ��D$P�L$<Ƅ$�   �S�����$�   PƄ$�   �^����L$<QP�D$|PƄ$�   �6����L$,QP�D$lPƄ$�   �������j j�PƄ$�   �w ���L$T��Ƅ$�   ������L$pƄ$�   �������$�   Ƅ$�   �����L$8Ƅ$�   ������r�L$�@Q�@Ƅ$�    �Ѓ��L$Ǆ$�   �����y�����t	V�_ ���Ƌ�$�   d�    Y^[�Ĩ   � V�t$���d! �����^� ���������Q� YË�`��`��`��` ��`$��`(��`,��`0��`4��`8��`<��`@�����������������������������4�A    �A    �A    �����V��~ �4u��r�v�@4� �Ѓ��F    �F    ^���������������̸   ����������̸   �����������3�� ������������ ������������̡�rV�@4��@$h�  �v���t$��r�t$�@4�t$�@�t$�v�Ѓ�2�^� ����������������t$��t$�t$�t$�P� ��������3�� ����������̸   � ��������� �������������Q��rU�@V�@ W�|$���3���=INIb�!  �  =SACbqt(=$'  t
=MicM�i  �E W���P$�   _��^]Y� �E �L$Q�L$Q�͉t$�t$�P��t�t$��r�t$�@4�u�@�Ѓ��   _��^]Y� =ARDb�  ��rS�@j ���   j���Ћء�rj �@j���   ���ЋL$����rj �@j���   �ЋL$��rj �@j���   ���t$�U PVWS���R[�   _��^]Y� �E ���P�   _��^]Y� =NIVb\tD=NPIbt-=ISIbuS�u ����  P���  P���V�   _��^]Y� �E W���P_^]Y� �E ���P�   _��^]Y� =cnyst	_��^]Y� ��rj �@hIicM���   ���ЋU WP���R _^]Y� ������������j�h�	d�    P��,V�`r3�P�D$4d�    ��~ ��   ��r�v�@4�@�Ѓ|$H t+��rP�F�I0�p�Al�Ѓ��L$4d�    Y^��8� ���L$ hARDb�D$�D$    �����NP�D$P�D$P�D$H    ��  ��r�L$���   Q� �Ѓ��L$ �D$<���������L$4d�    Y^��8� ����������̡�r�t$�@4�q�@l�Ѓ��   � ̡�r�q�@4�@�Ѓ�������������̡�r�q�@4�@�Ѓ�������������̡�r�q�@4�@�Ѓ�������������̡�r�q�@4�@|�Ѓ�������������̡�r�q�@4���   �Ѓ����������̡�r�t$�@4�q�@(�Ѓ�� �������t$��r�t$�@4�t$�@,�q�Ѓ�� ���������������t$��r�t$�@4�q�@0�Ѓ�� �̡�r�q�@4�@4��Y��������������̡�r�t$�@4�q���   �Ѓ�� ��̡�r�t$�@4�q�@ �Ѓ�� �����̡�r�t$�@4�q�@$�Ѓ�� �����̡�rV���   �t$�@WV���Ѓ�����rV���   u�@@�Ћ�rP�I4�w�A �Ѓ�_^� �@�Ѓ�����ru&���   V�@8�Ћ�rP�I4�w�A$�Ѓ�_^� �@h�3��0  h  �Ѓ�_^� ����������������t$��r�t$�@4�q�@D�Ѓ�� ���t$��r�t$�@4�q�@H�Ѓ�� ���t$��r�t$�@4�q�@L�Ѓ�� ���t$��r�t$�@4�q�@P�Ѓ�� �̡�rS���   V�@W�|$W���Ѓ�����r���   �@��   �t$V�Ѓ�����rV���   u5�@@�Ћ�rW���   ���I@�ы�rV�I4P�s�AP�Ѓ�_^[� �@�Ѓ�����ru<���   V�@8�Ћ�rW���   ���I@�ы�rV�I4P�s�AH�Ѓ�_^[� �@h�3��0  h�  �Ѓ�_^[� W�Ѓ�����r��   ���   �t$�@V�Ѓ�����rV���   u5�@@�Ћ�rW���   ���I8�ы�rV�I4P�s�AL�Ѓ�_^[� �@�Ѓ�����ru<���   V�@8�Ћ�rW���   ���I8�ы�rV�I4P�s�AD�Ѓ�_^[� �@h�3��0  h�  �Ѓ�_^[� �@h�3��0  h�  �Ѓ�_^[� ����������t$��r�t$�@0�t$���   �t$�q�Ѓ�� ��������t$��r�t$�@4�t$�@�t$�q�Ѓ�� �����������t$��r�t$�@4�t$�@�t$�q�Ѓ�� �����������t$(��r�t$(�@4�t$(�@T�t$(�t$(�t$(�t$(�t$(�t$(�t$(�q�Ѓ�,�( ���t$��r�t$�@4�t$��  �t$�q�Ѓ�� ������̡�rh�����@4h�����@Th�����t$�t$h����h����h����h�����t$(�q�Ѓ�,� ����������̡�r�t$�@4�q�@8�Ѓ�� �����̡�r�t$�@4�q�@<�Ѓ�� �������t$��r�t$�@4�q���   �Ѓ�� ��������������̡�r�q�@4�@@�Ѓ�������������̡�r�q�@4��  �Ѓ����������̡�r�D$�@4����  �$�q�Ѓ�� ����������t$��r�t$�@4�t$�@X�t$�q�Ѓ�� ���������̡�r�q�@4�@`��Y��������������̡�r�q�@4�@d�Ѓ���������������t$��r�t$�@4�t$��   �t$�q�Ѓ�� ��������t$��r�t$�@4�t$�@\�t$�t$�t$�q�Ѓ�� ���t$��r�t$�@4�q��  �Ѓ�� ����������������t$��r�t$�@4�q�@h�Ѓ�� ���t$��r�t$�@4�q��  �Ѓ�� ����������������t$��r�t$�@4�q�@p�Ѓ�� ��j�h
d�    P��VW�`r3�P�D$ d�    ��hYALf�L$����P��r�w�B4�D$0    �@l�Ѓ��L$�D$(���������L$ d�    Y_^�� ������������UVW�|$���t��r�L$�@j ���   j�Љ�t$��t��r�L$�@j ���   j�Љ��rV�@4W�u�@p�Ѓ�_^]� �������������t$��r�t$�I�@0�t$���   �q�Ѓ�� ���������t$��r�t$�@4�t$�@x�t$�q�Ѓ�� ���������̡�r�t$�@4�q�@t�Ѓ�� �������t$��r�t$�@4�t$���   �t$�t$�q�Ѓ�� ����t$��r�t$�@4�t$���   �t$�t$�q�Ѓ�� ��̃���rSW�D$    �D$    �@�ًL$$���   �{j j�ЋL$$�D$��rj �@j���   �ЉD$��r�L$�@0Q�@`�L$Q�w�С�r�s�@4�@�Ћ�rj �I0�T$,R�T$4R�T$(R�T$4RP�C�p�Ah�Ѓ�,�|$( _[t.�|$$ t.�L$�T$;�~C�D$�;�}9�$�T$;�~.�D$��|$$ u�L$�T$;�~�D$�;�}�   ��� 3���� ����������������t$�D$��r���@4�D$�D$���   �$�t$�q�Ѓ�� ������t$��r�t$�@4�t$���   �q�Ѓ�� ����������̡�r�q�@4���   �Ѓ�����������V��V�D4��rh�� �@0� �Ѓ��F�F    ��^�����V��N�D4��t��rQ�@0�@�Ѓ��F    ^������̸   ����������̸   ����������̸   � ��������3�� �����������3���������������� ����������������������������̡�rV�@W�|$�@ �����=NIVb��   ��   =TCAbttK=$'  t2=MicM��   ��rj �@hIicM���   ���ЋWP���R_^� �W���P_�   ^� ��rj �@hdiem���   ���ЋWP���R_^� =INIbuz�~ u���F   �P_^� �~ t�����P_^� =atni=t/=ckhct=ytsdu8����P_�F    3�^� ����P_^� �.�  _3�^� =cnys����_3�^� �����V��N��u3�^� ��rj �@0j ���   j j j �t$4j �t$(jQ���t$D��r�t$D�@0�t$D���   �t$Dj �t$D�v�Ѓ�D^� ��������̋I��u3�á�rQ�@0�@�Ѓ�����̋I��u3�� ��rQ�@0�@�Ѓ�� j�hW
d�    P��V�`r3�P�D$d�    �D$    �q��u �D$,�    �p�L$d�    Y^�� � �D$0�H���rQ�t$8�@0R���   �L$VQ�ЋЋt$@j �    �F    ��rR���   V�@�D$D   �Ћ�r�D$,���   P�	�D$,   �D$H �у�$�ƋL$d�    Y^�� � �������������̡�r�t$�@0�q���   �Ѓ�� ��̡�r�q�@0���   �Ѓ����������̡�rj �@0j ���   j j j j j j j4�q�Ѓ�(�������̡�rj �@0j ���   j j j j j j j;�q�Ѓ�(�������̡�r�t$�@0�q�@�Ѓ�� �����̋I��t(��rj �@0j ���   j j j j �t$j jQ�Ѓ�(� ���������������t$��r�t$�@4�t$�@,�q�Ѓ�� ���������������t$��r�t$�@4�q�@0�Ѓ�� �̡�r�q�@4�@4��Y���������������V�q��u3�^� �D$�H���rQ�t$�@0R�@V�Ѓ�^� ��������������V�q��u3�^� �D$�H���rQ�@0R���   V�Ѓ�^� ��������������̋D$3�h�����h  ���Pj BRj �t$ �t$ �   � ����j�h�
d�    P��$VW�`r3�P�D$0d�    ��htniv�L$ �k�����r�t$D�@hulav�@4�L$$�D$@    �С�rhgnlf�@htmrf�@4�L$$�С�r�t$H�@hinim�@4�L$$�С�r�t$L�@hixam�@4�L$$�С�r�t$P�@hpets�@4�L$$�С�r�t$T�@hsirt�@4�L$$�ЋL$X�t$\��  �u�����t.��rQ�@h2nim�@4�L$$�С�rV�@h2xam�@4�L$$�ЍD$P�t$D�D$P������P��r�D$<���   �@8�Ћ�r�����   �D$�	P�D$@ �у��L$�D$8�����d����ƋL$0d�    Y_^��0�  ��������������U����j�h�
d�    P��pV�`r3�P�D$xd�    ��htlfv�L$4�������r�E�@���@,�$hulav�L$<Ǆ$�       �С�r�u,�@htmrf�@4�L$8�С�r�E�@���@,�$hinim�L$<�С�r�E�@���@,�$hixam�L$<�С�r�E$�@���@,�$hpets�L$<�С�r�uD�@hsirt�@4�L$8���U0W�f.џ��Dz�E8f.����D{A��r���@�$�@,h2nim�L$<�С�r�E8�@���@,�$h2xam�L$<�С�r�u@�@hdauq�@4�L$8�ЍD$0P�u�D$$P������P��rƄ$�   ���   �@8�Ћ�r�����   �D$ �	PƄ$�    �у��L$0Ǆ$�   �����^����ƋL$xd�    Y^��]�@ ����������t$(W�j ���D$�$�D$8htemf�� �D$�D$T�D$�D$L�D$�D$D�$�t$@�����( �������L$f.05�5�% 5���D{�Y��^��T$f.85���D{�Y��^��t$(W�j ���D$�$�D$8�Y�hrgdf�� �^��D$�D$D�L$�T$�$�t$@�����( ���t$(�5W�j ���D$�$�D$8�^�htcpf�� �D$�D$T�^��D$�D$L�^��D$�D$D�$�t$@�����( ��U����j�h�
d�    P��hSVW�`r3�P�D$xd�    �ًE��u)��r�@���   �Ѕ�u�L$xd�    Y_^[��]� ���e  htlfv�L$4�������ufn�������YǄ$�       �D$�D$�$��s �F�\$$�D$�D$�$�s �D$$�\$�^D$��r�$�@hulav�@,�L$<�С�rhmrff�@htmrf�@4�L$8�Ћufn�������Y�D$$�D$$�$�Es �F�\$�D$$�D$$�$�*s �D$�\$$�^D$$��r�$�@hinim�@,�L$<�Ћufn�������Y�D$$�D$$�$��r �F�\$�D$$�D$$�$��r �\$$�D$�^D$$��r�$�@hixam�@,�L$<�С�r��2�@���@,�$hpets�L$<�С�rj �@hdauq�@4�L$8�С�rW�@hspff�@4�L$8�С�r�u �@hsirt�@4�L$8�ЍD$0P�u�D$$P������P��rƄ$�   ���   �@8�Ћ�r�����   �D$ �	PƄ$�    �у��L$0Ǆ$�   �����%����ƋL$xd�    Y_^[��]� ��������������j�hd�    P��$V�`r3�P�D$,d�    ��hCITb�L$������r�t$@�@hCITb�@8�L$ �D$<    �С�r�t$D�@hsirt�@4�L$ �С�r�t$H�@hulav�@4�L$ �ЍD$P�t$@�D$P���q���P��r�D$8���   �@8�Ћ�r�����   �D$�	P�D$< �у��L$�D$4���������ƋL$,d�    Y^��0� �����V�q��u3�^� �D$�D$�H���rQ�t$$�@0���@(�D$�D$(�$�t$$RV�Ѓ�$^� j�h&d�    P��V�`r3�P�D$d�    ��L$,�D$P�\���j �t$4��P�t$4�D$0    �b�����r���I�D$�IP�D$$�����у��ƋL$d�    Y^��� �������������V�q��u3�^� �D$�H���rQ�@0�L$�@,QRV�ЋL$3҃�9T$^�� ��������������V�q��u3�^� �D$�H���rQ�t$�@0R�@,V�Ѓ�^� ��������������V�q��u3�^� �D$�H���rQ�t$�@0R�@0V�Ѓ�^� ��������������UVW���O����   �D$�l$�P�0��rR�@0U�@0VQ�Ѓ���tb� t\�D$�H���rQ�p0�EP�F0R�w�Ѓ���t6���t/�D$�H���rQ�p0�EP�F0RW�Ѓ���t_^�   ]� _^3�]� �QV�q��u3�^Y� �D$W�H���rQ�L$�D$    �@0Q�@8RV�Ћ�����t=�T$��t5��r�t$�AR�@�Ћt$����t��rV�@�@��V�֥������_^Y� �����������V�q��u3�^� �D$�H���rQ�t$�@0�t$�@<RV�Ѓ�^� ���������̋D$��V���u��r�@���   �Ѕ�u^��� W���_^  �v����t#�D$$�H���rQ�@0�L$�@0QRV�Ѓ���fn�������Y(5�L$ �D$�D$�Y(5�$�.! �~ �L$,_f��~@��f�A^��� ��������������j�hId�    P��V�`r3�P�D$d�    ��r�L$�@Q�@�Ѓ��D$P�t$,���D$(    ��������t�L$,�D$P�I�����r�D$�IP�I�D$$�����у��ƋL$d�    Y^��� ������V�q��u3�^� �D$�H���rQ�@0j ���   j j j j j Rj1V�Ѓ�(^� ̡�rV�@j �t$���   ��L$��h���h  �j j jj P�t$$���%���^� ̡�rV�@j �t$���   ��L$���t$$���t$$j �t$(�t$(�t$(P�t$$�����^�  �������������U������<��rV�@�����   W��$�u��M���\$8�E8j �u@�΃��D$�E0�$�u,�E$�� �D$�E�D$�E�D$�D$t�$�u�����^��]�< ���������������U������<��rV�@�����   W��$�u��M���\$8j j ��W��D$�$�E$htemf�� ���D$�E�D$�E�D$�D$t�$�u�L���^��]�$ �����U������<��rV�@�����   W��$�u��M���\$8�Uf.05�5�% 5���D{�Y��^��Mf.85���D{�Y��^�j j ��W��D$�$�E$�Y�hrgdf�� ���^��D$�D$t�T$�L$�$�u�x���^��]�$ �U������<��rV�@�����   W��$�u��M���\$8�5j W�j �����D$�$�E$�^�htcpf�� �D$�E�^��D$�E�^��D$�D$t�$�u�����^��]�$ ̃�0��rV��W��D$��2�L$Q�t$H�D$�@�L$,���   Q�L$L���~ j �t$Tf�D$�t$T�~@�t$T�D$$P�t$P���t$Pf�D$8�����^��0� ���j�htd�    P�� V�`r3�P�D$(d�    ��r�L$�@Q�@�Ѓ��L$<�D$P�t$D�D$ P�D$<    �&K  �t$D��j P�t$D�D$@������r���I�D$�IP�D$4 �ѡ�r�L$�@Q�@�D$8�����Ѓ��ƋL$(d�    Y^��,� ���j�h�d�    P��HV�`r3�P�D$Pd�    ��L$4�Ѧ���L$dP�t$l�D$ P�D$d    ��I  �L$Q���D$\�U���j j P�t$l���D$h�`�����r���I�D$�IP�D$\�у��L$�D$X �U����L$4�D$X�����D����ƋL$Pd�    Y^��T� ���������������U������x�U��2V�uW���D$0���t.��r���@W����   �$R�����\$0�D$0�D$0��rW��L$8Q�u�D$@�D$H�D$P�@�L$p���   Q�����~ �wf�D$P�~@f�D$X�~@f�D$`��u
3�_^��]� �E�E�H���rQ�u �@0���@(�D$�D$H�$�L$hQRV�Ѓ�$_^��]� ���V�q3���t,�D$�H���rQ�@0�L$�@,QRV�Ћ�3���9D$����rP�Q�t$�L$�R0�ҋ�^� �������������V�q��t#�D$�H���rQ�@0�L$�@,QRV�Ѓ�����r�t$�A�t$�L$�@4�Ћ�^� ����̃�V�q��t#�D$�H���rQ�@0�L$�@0QRV�Ѓ�����r�D$�A�L$�@,���$�t$ �Ћ�^��� ����̃�V�D$P�t$ W��t$ �D$��2�D$�������r���Q�L$ �R@�D$P�t$(�ҋ�^��� ������������̃�V��W�~W��D$�D$�D$����   �D$$�H���rQ�@0�L$�@0QRW�Ѓ���t�~��tx�D$(�H���rQ�@0�L$�@0QRW�Ѓ���tS�v��tL�D$,�H���rQ�@0�L$�@0QRV�Ѓ���t'��r�L$�@Q�t$8�L$8�@H��_�   ^��� _3�^��� �����������j�h�d�    P��V�`r3�P�D$d�    ��r�L$�@Q�@�Ѓ��D$P�t$,���D$(    ������r���Q�L$,�R8�D$P�t$4�ҡ�r�L$�@Q�@�D$$�����Ѓ��ƋL$d�    Y^��� ��������������j�h�d�    P��V�`r3�P�D$$d�    ��L$�����D$P�t$8���D$4    ������r���Q�L$8�R<�D$P�t$@�ҍL$�D$,����諣���ƋL$$d�    Y^��(� �����̃� V�qW��D$�D$�D$��t(�D$(�H���rQ�@0�L$�@<Q�L$QRV�Ѓ����T$0���t��r�A�L$�@HQ�L$0R�ЋT$4���t ��r�D$�@�L$,�@,���$R�Ћ�^�� � ����̋D$3҃8V�p�¸   h���h  ���E�3�����Rj @Pj V�t$$����^� �T$�t$3��:�t$��P�t$ �t$ �t$ �r�t$ ����� �T$�D$03��:��P�t$<���D$�D$@�$�t$<�D$8�� �D$�D$P�D$�D$H�D$�B�$�t$@�����8 ���̋D$3҃8�H��W�Rj ���D$�$�D$4htemf�� �D$�D$P�D$�D$H�D$�$�t$@�Q����  �������������̋D$�T$�h�5�% 53҃8��f.05���D{�Y��^��L$f.85���D{�Y��^�Rj ��W��D$�$�D$4�Y�hrgdf�� �^��D$�T$�L$�,$�t$@�����  ���������̋D$�53҃8W����PRj ���D$�$�D$4�^�htcpf�� �D$�D$P�^��D$�D$H�^��D$�$�t$@�����  ���������̋T$3��:��P�t$�B�t$�t$P�t$�t$�V���� ��̋D$�t$3҃8��RP�t$����� ���������������j�h(d�    P��$V�`r3�P�D$,d�    ��hgnrs�L$�|����D$@�D$4    �D$   �D$��r�L$�@Q���   j�L$ �D$<�С�r�L$���   Q� �D$8 �ЋD$H���D$   �D$��r�L$�@Q���   j�L$ �D$<�С�r�L$���   Q� �D$8 �Ѓ��D$P�t$@�D$P������P��r�D$8���   �@8�Ћ�r�����   �D$�	P�D$< �у��L$�D$4����������ƋL$,d�    Y^��0� �����������W�y��u3�_� �D$�D$�H���rV�p0�D$Q�t$(�����D$�D$,�$P�F(RW�Ѓ�$^_� ���������̡�rj �@0j ���   j j j j j j j �q�Ѓ�(�������̋I��u3�� ��r�t$�@4�t$��  Q�Ѓ�� ����̋I��u3�� ��r�t$�@4�t$�@hQ�Ѓ�� �������̋I��u3�� ��r�t$�@4�t$�@pQ�Ѓ�� �������̋I��u3�� ��r�t$�@4�t$��  Q�Ѓ�� ������t$��r�t$�@0�t$���   �t$�q�Ѓ�� ������̡�r�P0�D$�pj j j �t$�t$j �0���   j=�q�Ѓ�(� �����������̡�r�P0�D$�p�t$j j j��t$j �0���   j=�q�Ѓ�(� �����������̋D$�t$���|rEС�r�2�@0�t$�@@�q�Ѓ�� ��Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$jQ�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$jQ�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj �t$$�D$    �t$ �@0�t$ ���   �t$ �t$0�t$$jQ�ЋD$(��(Y� ��������������Q�I��u3�Y� ��r�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j*Q�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� ��Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� ��Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$j	Q�ЋD$(��(Y� ��Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$j
Q�ЋD$(��(Y� ��Q�I��u3�Y� ��r�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$j'Q�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   �t$0�t$$j,Q�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j:Q�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj j j �t$�D$    �t$ �@0j ���   j j)Q�ЋD$(��(Y� ������Q�I��u3�Y� ��r�$Rj j �t$�D$    �@0j �t$ ���   j j j)Q�ЋD$(��(Y� �����̋I��u3�� ��rj �@0j ���   j �t$�t$�t$j �t$ jQ�Ѓ�(� ���Q�I��u3�Y� ��r�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$jQ�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj �t$ �D$    �t$ �@0�t$ ���   �t$ j �t$$j>Q�ЋD$(��(Y� Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� �̡�rj �@0j ���   j �t$�t$�t$j �t$ j.�q�Ѓ�(� �������������V�q��u3�^� �D$�H���rQ�@0j ���   j j j �t$ �t$(RjV�Ѓ�(^� �������������V�q��u3�^� �D$�H���rQ�@0j ���   j j j j j RjV�Ѓ�(^� �V�q��u3�^� �D$�H���rQ�t$�@0R�@\V�Ѓ�^� �������������̃�SVW�t$ �ٍL$�+
 �D$ P�D$P�L$�h
 ��tm�|$�L$ ��tJ��rQ���   �@H�ЋS������tR�w��rj �A0j ���   j j �t$ V�7jR�Ѓ�(��t%�D$ P�D$P�L$��	 ��u�_^�   [��� _^3�[��� ��������������Q�I��u3�Y� ��r�$Rj j �t$ �D$    �t$ �@0�t$ ���   j �t$$jQ�ЋD$(��(Y� �̡�rV�@4W�|$� �w���ЋD$�G    �w�H���rQ�t$�@0W���   R�v�Ѓ�3Ʌ����G_^��� �������̋I��u3�� ��rj �@0j ���   j �t$�t$�t$j �t$ j/Q�Ѓ�(� ��̋T$��u3�� �r�B    ��r�t$�@0�q���   �Ѓ�� �����������̋I��u3�� ��rj �@0j ���   j j j �t$j j jQ�Ѓ�(� ��������̡�rj �@0j ���   j j j j j j j6�q�Ѓ�(�������̋I��u3�� �t$��r�t$�@0�t$�@DQ�Ѓ�� ���̋I��u3�� �t$��r�t$�@0�t$�@H�t$�t$�t$Q�Ѓ�� �������̋I��u3�á�rQ�@0�@X�Ѓ�����̋I��u3�� ��r�t$�@0�t$�@LQ�Ѓ�� �������̋Q��u3�� ��r�H0�D$   �P�APR�Ѓ�� �����̋I��u3�� ��r�t$�@0Q�@P�Ѓ�� �����������̋I��u3�� �t$��r�t$�@0�t$�@T�t$Q�Ѓ�� j�hKd�    P��VW�`r3�P�D$ d�    ���L$萳���D$0�L$�P�0��rR�@0Q���   j j j j j Vj8�w�D$P    �Ћ���(��t�L$4�D$P貳���L$�D$(����葳���ƋL$ d�    Y_^�� � ����������̋D$V�P�0��rR�t$�@0j ���   j j j j Vj9�q�Ѓ�(^� ���������̋D$V�P�0��rR�t$�@0�t$�@h�t$�t$V�q�Ѓ�^� �������������UVW�|$���t��r�L$�@j ���   j�Љ�t$��t��r�L$�@j ���   j�Љ��rV�@0W�u�@`�Ѓ�_^]� �������������t$��r�t$�@0�t$���   �q�Ѓ�� ����������̋T$��r�@0��t*���   R�q�Ћ�r�t$�ЋA0R���   �Ѓ�� �t$�@|�q�Ѓ�� �����t$��r�t$�@0�t$�@p�t$�t$�q�Ѓ�� �������t$��r�t$�@0�t$�@d�t$�t$�q�Ѓ�� �����̡�rj �@0j �t$���   �t$ �t$ �t$j �t$ j3�q�Ѓ�(� ����������̋D$j ���rj �@0j ���   j j j j Rj�q�Ѓ�(� �D$j ���rj �@0j ���   j j jj Rj�q�Ѓ�(� �D$j ���rj �@0j ���   j j j j Rj�q�Ѓ�(� �D$V�P�0��rR�@0j ���   j j j j j Vj"�q�Ѓ�(^� �����������̋D$V�P�0��rR�@0j ���   j j j j j Vj5�q�Ѓ�(^� �����������̋D$V�P�0��rR�@0j ���   j j j �t$ j Vj<�q�Ѓ�(^� ���������̡�rV�@0j ���   j j j j �t$ ��j �t$$j�v�С�r�t$8�@0�v�@t�Ѓ�0^� ��������̡�rj �@0j ���   j j j j j j j�q�Ѓ�(�������̡�rj �@0j ���   j j j j �t$j j�q�Ѓ�(� ��̡�rj �@0j ���   j j j j j j j�q�Ѓ�(�������̡�rj �@0j ���   j j j j j �t$ j�q�Ѓ�(� ��̡�rj �@0j ���   j j j j �t$ �t$ j&�q�Ѓ�(� ̡�rj �@0j ���   j j j j j j j(�q�Ѓ�(�������̡�rj �@0j ���   j j j j j j j#�q�Ѓ�(�������̡�rj �@0j ���   j j �t$�t$j �t$ j+�q�Ѓ�(� ��������������̡�rj �@0j ���   j j j j j j j0�q�Ѓ�(�������̡�r�t$�@0�q���   �Ѓ�� ���j�hnd�    P��V�`r3�P�D$d�    ���t$D�L$荭����r�t$0�@h8kds�@4�L$�D$,    �С�r�L$DQ�L$Qj �t$L�D$T    �t$L�@0�t$L���   �t$L�t$Hj2�v�Ћt$l��(�L$�D$$�����6����ƋL$d�    Y^�� � ̡�r�q�@0���   �Ѓ����������̋I��u3�� ��rj �@0j ���   j j j j j �t$ j-Q�Ѓ�(� ��������̃���rW�@j ���   ���L$(j�ЋL$$�D$��rj �@j���   �ЉD$��r�L$�@0Q�@`�L$Q�w�С�r�T$�H0�D$,�pR�T$,R�T$$R�T$0R�0�Ah�w�Ѓ�(�|$( _t.�|$( t.�L$�T$;�~C�D$�;�}9�$�T$;�~.�D$��|$( u�L$�T$;�~�D$�;�}�   ��� 3���� ��SV�t$W��u�q��r�\$�@j ���   hdiuM���Ћ���tH;>u_^3�[� ��rj �@hIicM���   ����;�u��rj �@h1icM���   ���Шu��>_^�   [� ������������j�h�d�    P��V�`r3�P�D$d�    ��r�t$,�@hfnic�@T���ЋЅ�t��rj
�A�ʋ��   �Ѕ���   hfnic�D$P���(  �t$0P���D$(    �̪���L$�D$$����諪����r�΋@�@ �Ѓ��t��r�΋@�@ �Ѕ�u��rhfnic�@�΋@$�С�r�t$4�@j
�@8���ЋL$d�    Y^�� ����������̡�r�q�@0���   �Ѓ�����������j�h�d�    P��$V�`r3�P�D$,d�    ��hmnrs�L$謩����r�t$@�@j�@4�L$ �D$<    �ЍD$P�t$@�D$P�������P��r�D$8���   �@8�Ћ�r�����   �D$�	P�D$< �у��L$�D$4�����q����ƋL$,d�    Y^��0� ������������j�h�d�    P��$V�`r3�P�D$,d�    ��|$@ �SSSS�DSSSE�P�L$�Ψ����r�L$�@�D$4    �@ �Ћ�rj�QP�B4�L$ �ЍD$P�t$@�D$P�������P��r�D$8���   �@8�Ћ�r�����   �D$�	P�D$< �у��L$�D$4����脨���ƋL$,d�    Y^��0� ���������������V��V�D4��rh�� �@0� �Ѓ��F�F    �l4�F   �F    ��^�V��N�D4��t��rQ�@0�@�Ѓ��F    ^�������V��N�F    ��tk��rj �@0j ���   j j j j j j jQ�С�r�t$<�H0�t$<3�9D$H�t$<���t$<j ��
P�v���   �Ѓ�D��t�~ t	�   ^� 3�^� �������������̋D$�A�I��u3�� ��rQ�@0�@�Ѓ�� ��������̡�rS�@�\$�@ V�����=ckhc��   tz=cksata=TCAb��   ��rW�@j ���   hdiem���Ћ��SW���F   �R�~ ��t��t��u3�������P�L���_^��[� �~ tg����P^[� �~ tU��rj �@0j ���   j j j j j j j �v�Ѓ�(��t)�F    ^�   [� =atnit�t$��S�l���^[� ^3�[� U��} ��   S�\$V�t$W�|$$��wy�$�� 9t$��   �f9t$��   �Z9t$��   �N9t$��   �B�D$;�~:;���   �0�D$;�|(;�~~�"�D$;�|;�|p��D$;�~;�~b�9t$uZ��rj �@0j ���   j j j j j �t$0j�u��fn������(j���D$fn�����$S�6W  ���E    _^[]� �� $� 0� <� H� Z� h� v� �� W��� �\  V�t$����   �$��� �D$f/D$�4  ��   �D$f/D$�  ��   �L$f/L$�  �   �L$f/L$��   �   �T$f/T$��   �D$$f/���   �n�T$f/T$r`�D$$f/���   �N�T$f/T$r@�D$$f/���   �.�T$f/T$v �D$$f/�sl��D$f.D$���DzX��rj �@0j ���   j j j j j �t$(j�w���D$L��(�t$,���D$�D$0�$V�U  ���G    ^_�$ �I 2� I� `� w� �� �� Һ � � �������������D$j���D$�D$0�D$�D$(�$�t$$�t$$�+����  ���������D$j���D$�D$0�D$�D$(�$�t$$�t$$������  ���������D$j���D$�D$0�D$�D$(�$�t$$�t$$�����  ��������V��V�D4��rh�� �@0� �Ѓ��F�F    ��4�F   ��^��������V��N�D4��t��rQ�@0�@�Ѓ��F    ^������̡�rV�@��L$�@ ��=cksat]=ckhct�t$���t$�?���^� j j j j j j �F   ��rj �@0j ���   j �v�Ѓ�(��t!�F    �   ^� �~ t����P^� 3�^� �j�h
d�    PQV�`r3�P�D$d�    ��t$�D4��rV�@0h�� � �Ѓ��F�F    �F   �D$ �L$��4�F��rj �@hmyal���   �D$    �ЉF��t��t�F    ��r�L$�@j
���   hhfed�ЉF�ƋL$d�    Y^��� ����̡�rV�@��L$�@ ��=ytsdt�t$���t$�v���^� ��r�v�@0���   �Ћ�����P�   ^� ������������3���������������3�������������������������������3���������������3���������������3���������������3�� �����������Q�L$�$    �?  �D$Y� ������̋A��uË ���������������������V���PD��t�D$9Ft
�F����PH^� ������������̋A�������������j0�t$�uK  ����j0�t$�e�  ��P�\K  �����������j�h-d�    P���`r3�P�D$d�    �t$(�D$�t$(P�K�  j0P�D$0    �K  ��r�L$�@Q�@�D$4�����Ѓ��L$d�    Y�����������������j�hPd�    P���`r3�P�D$d�    �t$,�D$�t$,�t$,P藓  j0P�D$4    �J  ��r�L$�@Q�@�D$8�����Ѓ��L$d�    Y�������������j$�t$�EJ  3Ƀ���������������j$�t$�%�  ��P�J  3Ƀ����������������������j�hsd�    P��S�`r3�P�D$d�    �t$,�D$�t$,P���  j$P�D$4    �I  ��r3ۋI���I�D$P���D$8�����у��ËL$d�    Y[����j�h�d�    P��S�`r3�P�D$d�    �t$0�D$�t$0�t$0P�F�  j$P�D$8    �6I  ��r3ۋI���I�D$ P���D$<�����у��ËL$d�    Y[���������������̡�r�t$�@�t$���   j �Ѓ�����t$��r�t$�@�t$���   j �Ѓ���������������̡�r�@���  �࡜r�@0���   ��j�h�d�    P��VW�`r3�P�D$ d�    �t$8�D$    ��r�t$8�@0�L$���   Q�Ћ���r�|$<�IW�I�D$8   �ѡ�rW�@V�@�Ћ�r�D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� ����j�hd�    P��(SUVW�`r3�P�D$<d�    �D$    ��r�|$L�@W�@�D$H    �Ѓ���r�L$P�@3ۋ��   SS�D$L    �D$    �ЋL$P�D$��rS�@j���   �Ћ����&  3���I ��~|��r�L$�@Q�@�С�rj �@j��@�L$(h4Q�Ѓ���r�ϋ@�D$D   �@<�Ћȡ�rj��@j��@L�T$$RQ���С�r�L$�@Q�@�D$H �Ѓ�V�t$�D$4P�!�������r�ϋ@�D$D   �@<�Ћȡ�rj��@j��@LVQ���С�r�L$,�@Q�@�D$H �С�r�L$T�@�����   j ��
UC�ЉD$��rj �P�M���   Q�L$X�ҋ���������ǋL$<d�    Y_^][��4�����������̡�r�@0���   �࡜r�@0���   �࡜r�@0���   ����W��JR��A(�P$j j h����I  �������������̸3�����������j�had�    P��8SVW�`r3�P�D$Hd�    ����L$Q���P(���W�D$P    ��t&��rj �A0j ���   j j j j Vj jR�Ѓ�(��r�L$�@Q�@�D$T�����С�r�L$�@Q�@�Ѓ��O�D$P   ��t ��rj �@0�T$�@HRj jj?j Q�Ѓ���r�L$�@Q�@�D$T�����С�r�L$�@Q�@�Ѓ��O�D$P   ��u3��>��r�T$Rj j j h  
 j�T$,R�D$,    �@0h�  ���   jQ�ЋD$8��(����r�L$�@Q�@���D$T�����Ѓ���t3��L$Hd�    Y_^[��Dá�r�L$�@Q�@�Ѓ��O�D$P   ��t ��rj �@0�T$�@HRj j j8j Q�Ѓ���r�L$�@Q�@�D$T�����ЋO����t��rj�@0Q�@P�Ѓ��L$4�(�������r�D$$�IP�I�D$T   �у�Vh   h  K j;�D$4Ph	��h�  ���D$l�`�����r�L$$�@Q�@�D$T�Ѓ��L$4�D$P���������O��t��rQ�@0�@X�Ѓ��O��t��rQ�@0�@X�Ѓ��O��t&��rj �@0j ���   j j j jj j jQ�Ѓ�(j�$��A  ���   �L$Hd�    Y_^[��D����j�h�d�    P��VW�`r3�P�D$$d�    ��j�N��  �F4    �F8    �F<    W��F(��rh�   �@0�v�@�С�r�L$�@Q�@�С�rj �@j��@�L$(h$3Q�Ѓ�j j �D$P�D$P���D$<    �D$�  �D$     �п����r�L$�@Q�@�D$0�����Ѓ��Nj j�'�  �L$$d�    Y_^��$������j�h�d�    P��\VW�`r3�P�D$hd�    ��r�L$�@Q�@�С�rj �@j��@�L$ hh3Q���F(�Y5Ǆ$�       �D$ �  �D$$    �,�P�D$LP��Y���L$0QP�D$HPƄ$�   �  ��(j j P�D$P��Ƅ$�   �Ѿ����r�L$$�@Q�@�D$t�С�r�L$8�@Q�@�D$x �С�r�L$�@Q�@�D$|�����Ѓ��L$Thtats�8�����rj�@j�@0�L$\�D$x   �С�r�F(�@�@,���L$\�$j�ЍD$TP�D$P�D$LP���D$�  �D$    �%�����r�L$D���   Q� �Ѓ��~4 t_��r�N0�@P�@h�ЋF4��t�v8�Ѓ��F<�F8    �F4    ���rhl3�@h�  ��0  �Ѓ���r�N0�@P�@l�ЍL$T�D$p����舓���L$hd�    Y_^��h� ����j�h�d�    P��@VW�`r3�P�D$Ld�    ����r�t$\�@�΋@ ��=MicMtg=fnic�  j�L$<�ْ���L$`P�D$X    �����L$8�D$T�����������r�L$`�@j�@4j�и   �L$Ld�    Y_^��L� ��rj �@hIicM���   ����=�����   htats�L$(�V�����rj �@j�@0�L$,�D$\   �ЍD$$P�D$P�D$P���D$�  �D$    �c�����r�L$���   Q� �Ѓ��L$$�D$T�����+����O�G   ��t��rQ�@0�@�Ѓ��t$`��V������L$Ld�    Y_^��L� �����������̃l$V��t3�^� j�N�v�  j��<  �N���F    ��t��rQ�@0�@�Ѓ��   ^� ����j���6�  j�<  ��3������������D$�A(� �̍A�������������VW��~4 tC��    ��rh(3�@hs  ��0  ��j
�OG  ��r�v �@P�@�Ѓ���uM9F4uá�r�N0�@P�@h�Ѓ~4 t9��rhH3�@h�  ��0  �С�r���@P�N0�@l���o���_3�^� �D$�F8�D$�F4��rS�@P�N0�@l�Ѓ~4 t#j
�F  ��r�v �@P�@�Ѓ���u89F4uݡ�r�N0�@P�@h�Ћ~<�F<    ��r�N0�RP�Rl��[��_^� [_3�^� �j�hd�    P��V�`r3�P�D$d�    �L$裏���L$0��r�D$$    ��t"�@4Q�@�Ѓ���t'��L$Q�t$8���R(�'�@0�t$,�@�Ћȃ���u3��?��T$R�t$8�P ��r�L$�@�@ �Ѓ��t��r�L$�@0Q�t$0�@x�Ѓ��L$�D$$�����c����ƋL$d�    Y^�� á�rV�@j �t$���   ��L$�Ћ���u�    �F^� ��u9Ft�   ^� ������������V�t$W��;t$u��r�L$�@j ���   htsem�Ѕ�u`��r�L$�@j ���   hrdem�Ѕ�uA�D$�D$�H��t2��rj �@0�T$�@,RVQ�Ѓ���t�t$���m
  _�   ^� _3�^� ������������j�h@d�    P��0VW�`r3�P�D$<d�    ����r�L$�@Q�@�С�r�L$ �@Q�@�D$L    �Ѓ��L$L�D$P�t$T�D$4P�D$P��  �Ћ�r�D$D�A�L$�@QR�С�r�L$4�@Q�@�D$P�С�r�L$(�@Q�@�D$T �С�r��@V�@�С�r�L$ �@V�@Q�Ѓ����
  ��r�L$�@Q�@�D$H�����Ѓ��L$<d�    Y_^��<� �������j�hcd�    P��SV�`r3�P�D$$d�    �ًt$<;t$@��   ��r�L$8�@j ���   htsem�Ѕ���   ��r�L$8�@j ���   hrdem�Ѕ���   ��r�L$�@Q�@�Ѓ��L$4�D$P�D$P�D$4    �t$�D$    �ٹ����u3��5��r���@��@V�С�r�L$(�@V�@Q�Ѓ����	  �   ��r�D$�IP�I�D$0�����у��ƋL$$d�    Y^[��$� 3��L$$d�    Y^[��$� �̡�rV�@j �t$���   ��L$�Ћ���u�    �F^� ��u9Ft�   ^� �����������̃�V�t$W��;t$ uy��r�L$�@j ���   htsem�Ѕ�uZ��r�L$�@j ���   hrdem�Ѕ�u;�L$�D$�D$�D$P�D$P�t$�"�����t�t$���#  _�   ^��� _3�^��� �����������̃���rV�@�����   W��$�t$��L$���\$����u�D$�    �F^��� ��u�Ff.D$���D{�   ^��� �̃�SV�t$��;t$ ��   ��r�L$�@j ���   htsem�Ѕ�ur��r�L$�@j ���   hrdem�Ѕ�uS�D$W��H�D$��t?��rj �@0�T$�@0RVQ�Ѓ���t"�D$�����$�'  ^�   [��� ^3�[��� ��0��rV��W��L$Q�t$@�D$�D$�D$�@�L$$���   Q�L$D���~�~P�~H����uf�^f�V�    f�N^��0� ��u3�Ff.ß��Dz�Ff.��Dz�Ff.����D{�   ^��0� ���̃�4�D$@S�\$HV�t$TW�|$T�L$;�t;�t;���   ��r�L$H�@j ���   htsem�Ѕ���   ��r�L$H�@j ���   hrdem�Ѕ���   �L$D�D$�D$�D$$�D$(P�D$P�D$ PW��D$,P�D$8�D$@�D$H�t$ �|$(�\$0�6�����t<�~D$(�L$����f� �~D$Hf�@�~D$Pf�@�  �   _^[��4� _^3�[��4� ����������̃�0��rV��W��D$��2�L$Q�t$@�D$�@�L$,���   Q�L$D���~ �~H�f�D$f�L$���uf�F�    f�N^��0� ��u�D$P�FP�  ����t�   ^��0� �������̃�SV�t$0��;t$4��   ��r�L$(�@j ���   htsem�Ѕ���   ��r�L$(�@j ���   hrdem�Ѕ�uh�L$$�D$�D$P�t$0W��D$��2�D$P�D$$�t$�#�����t.�~D$���ċ�f� �~D$(f�@�  �   ^[��� ^3�[��� �������j�h�d�    P��V�`r3�P�D$d�    ��t$�V�    �B    �D$$    ������D$    �D$    ��rj ���   �L$�@QR�D$0�С�r�L$���   Q� �D$4 �Ѓ��ƋL$d�    Y^�� ������������̡�rQ���   � ��Y��������������̃�V�t$W�|$ �f.���Dz�Ff.G���D{a�G�Y����D$�D$�$�E! �F�\$�Y�D$�D$�$�&! �D$�\$��f.D$���D{_�   ^���_3�^���������������j�h�d�    PQV�`r3�P�D$d�    �D$    ��r�t$�@V�@�D$    �С�rV�@�t$(�@�Ѓ���r�΋@�D$    �@<�D$   �Ћ�rj��Qj��t$,�RLP���ҋƋL$d�    Y^���������������V��N�D4��t��rQ�@0�@�Ѓ��D$�F    t	V�X������^� ��V��~ �4u��r�v�@4� �Ѓ��D$�F    �F    t	V��W������^� ����������̋���u�D$�    �A� ��u�A;D$t�   � ��̋���u�D$�    �A� ��u�Af.D$���D{�   � ������̋���u*�~D$f�A�~D$f�A�~D$�    f�A� ��u9�Af.D$���Dz"�Af.D$���Dz�Af.D$���D{�   � ���������������V�����u �~D$f�F�~D$�    f�F^� ��u�D$P�FP���������t�   ^� ���j�h�d�    PV�`r3�P�D$d�    ���D$    ���u!�    ��r�N�@Q�@�L$Q�Ѓ��#��u��r�T$�@�N�@xR�Ѕ�t�   ��r�L$�@Q�@�D$�����Ѓ��L$d�    Y^��� ����������j�hAd�    P���`r3�P�D$d�    �t$0�D$    ��r�T$�@R�@P�ЋL$,P�D$(   譁���L$�D$   �D$$ 跁���D$,�L$d�    Y��$� �j�h�d�    P�� �`r3�P�D$$d�    �t$<�D$    ��r�t$<�@�T$���   R�ЋL$4P�D$0   ��]���L$�D$   �D$, �P^���D$4�L$$d�    Y��,� ����������j�h�d�    P��VW�`r3�P�D$ d�    �t$8�D$    ��r�t$8�@�T$���   R�Ћ���r�|$0�IW�I�D$,   �ѡ�rW�@V�@�Ћ�r�D$�IP�I�D$   �D$8 �у��ǋL$ d�    Y_^�� � ̡�rQ�@L���   �Ѓ������������̡�r�t$�@L�t$���   Q�Ѓ�� ̡�rV�@L�񋀠   V�Ћȡ�r����u�@LQ�t$���   V�Ѓ�^� ���   �@P�Ћ�rP���   �L$�BH��^� ̡�rQ�@L��(  �Ѓ������������̡�r�t$�@L�t$��,  Q�Ѓ�� ̡�r�@L� �����̡�rV�@@�t$�@�6�Ѓ��    ^�̡�r�@L���   �࡜rV�@@�t$�@�6�Ѓ��    ^��j�h�d�    P���`r3�P�D$d�    �t$0�D$    ��rQ�@L�L$�@Q�Ѓ��L$,P�D$(   �~���L$�D$   �D$$ �~���D$,�L$d�    Y��$� ������������̡�r�t$�@L�t$�@Q�Ѓ�� ���̡�r�t$�@LQ���   �Ѓ�� ����̡�rQ�@L�@�Ѓ���������������̡�rQ�@L�@�Ѓ���������������̡�rQ�@L�@�Ѓ�����������������t$��r�t$�@L�t$�@ Q�Ѓ�� ��r�t$�@LQ��4  �Ѓ�� ������t$��r�t$�@L�t$�@$Q�Ѓ�� �t$��r�t$�@L�t$�@(�t$Q�Ѓ�� �����������̡�rQ�@L�@,�Ѓ���������������̡�rQ�@L�@0�Ѓ���������������̡�rQ�@L�@4�Ѓ���������������̡�rj �@LQ�@8�Ѓ�������������̡�r�t$�@L�t$��  Q�Ѓ�� ̡�r�@L���   �࡜r�@L���   �࡜r�@L��l  �࡜r�@L���   �࡜r�@L���   �࡜r�@L���   �࡜r�@L���   �࡜r�@L���   �࡜r�@L���   �࡜r�t$�@LQ�@<�Ѓ�� �������̡�r�@L���   �࡜rQ�@L�@��Yá�r�t$�@L�t$�@@Q�Ѓ�� ���̡�rj �@L�t$�@DQ�Ѓ�� �����̡�rj�@L�t$�@DQ�Ѓ�� �����̡�rj �@L�t$�@HQ�Ѓ�� �����̡�rj�@L�t$�@HQ�Ѓ�� �����̡�rQ�@L���   �Ѓ�������������j�h5d�    P���`r3�P�D$d�    �t$0�D$    ��rQ�@L�L$��  Q�Ѓ��L$,P�D$(   �z���L$�D$   �D$$ ��z���D$,�L$d�    Y��$� ����������j�h`d�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �[�  j �D$$P�D$P���D$D�C|�����L$���D$8 ���  ��t3����r�L$ ���   Q�@8�Ѓ�����r�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h�d�    P��$V�`r3�P�D$,d�    ���D$   �D$$   �D$P�L$�D$8    �D$�  �D$    �D$    �l  j�D$ P�D$P���D$@�d{���L$�D$4 �ր  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0�������j�h�d�    P��(SV�`r3�P�D$4d�    ���D$    �D$$    �D$,    �D$P�L$�D$@   �D$�  �D$     �D$$    �~  j �D$(P�D$P���D$H�z�����L$���D$<��  ��t�L$D�{S���"��r�L$$���   Q�@L�ЋL$H��P��T����r�D$$���   P�	�D$   �D$@ �ыD$H���L$4d�    Y^[��4� ����������j�hd�    P��(SV�`r3�P�D$4d�    ���D$    �D$$    �D$,    �D$P�L$�D$@   �D$�  �D$     �D$$    �}  j �D$(P�D$P���D$H�{y�����L$���D$<��~  ��t�L$D�kR���"��r�L$$���   Q�@L�ЋL$H��P�S����r�D$$���   P�	�D$   �D$@ �ыD$H���L$4d�    Y^[��4� ����������j�h>d�    P��$V�`r3�P�D$,d�    ��r�t$<�D$     �D$(    ���   �L$ �@(Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �p|  j�D$ P�D$P���D$@�hx���L$�D$4 ��}  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�hid�    P��$V�`r3�P�D$,d�    ��r�t$<�D$     �D$(    ���   �L$ �@(Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �{  j�D$ P�D$P���D$@�w���L$�D$4 ��|  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h�d�    P��,SV�`r3�P�D$8d�    ���D$(    �D$0    �D$P�L$�D$D    �D$ �  �D$$    �D$(    ��z  j �D$,P�D$P���D$L�v�����L$���D$@ �0|  ��tW��D$�D$���r�L$(���   Q�@<�Ѓ���r�\$�L$(���   Q� �D$D�������D$���L$8d�    Y^[��8�������������j�h�d�    P��V�`r3�P�D$$d�    ���D$4�D$   �D$�D$P�L$8�D$0    �D$�  �D$    �D$    ��y  j�D$P�D$<P���D$8��u���L$4�D$, �2{  ��r�L$���   Q� �D$0�����Ѓ��L$$d�    Y^��(� j�h�d�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �y  j �D$$P�D$P���D$D��t�����L$���D$8 �pz  ��t3����r�L$ ���   Q�@8�Ѓ�����r�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�hd�    P��$V�`r3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    �x  j�D$ P�D$P���D$@�t���L$�D$4 �y  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�h@d�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �[w  j �D$$P�D$P���D$D�Cs�����L$���D$8 ��x  ��t:��r�t$@���   W��	���2�D$ P�F�D$<�����у��K��r�L$ ���   Q�@P���~ �t$D��rf��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�hkd�    P��$V�`r3�P�D$,d�    ��r�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �v  j�D$ P�D$P���D$@�r���L$�D$4 �zw  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h�d�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �Ku  j �D$$P�D$P���D$D�3q�����L$���D$8 �v  ��t:��r�t$@���   W��	���2�D$ P�F�D$<�����у��K��r�L$ ���   Q�@P���~ �t$D��rf��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�h�d�    P��$V�`r3�P�D$,d�    ��r�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    � t  j�D$ P�D$P���D$@��o���L$�D$4 �ju  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� �������̡�r���@Lj�t$���   Q�L$Q�ЋL$$�~ f��~@f�A���� � ��̡�r���@Lj �t$���   Q�L$Q�ЋL$$�~ f��~@f�A���� � ���j�h�d�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �r  j �D$$P�D$P���D$D�n�����L$���D$8 � t  ��t:��r�t$@���   W��	���2�D$ P�F�D$<�����у��K��r�L$ ���   Q�@P���~ �t$D��rf��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�hd�    P��$V�`r3�P�D$,d�    ��r�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �pq  j�D$ P�D$P���D$@�hm���L$�D$4 ��r  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�hBd�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �p  j �D$$P�D$P���D$D�l�����L$���D$8 �r  ��t:��r�t$@���   W��	���2�D$ P�F�D$<�����у��K��r�L$ ���   Q�@P���~ �t$D��rf��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�hmd�    P��$V�`r3�P�D$,d�    ��r�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �`o  j�D$ P�D$P���D$@�Xk���L$�D$4 ��p  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�h�d�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �n  j �D$$P�D$P���D$D�j�����L$���D$8 � p  ��t3����r�L$ ���   Q�@8�Ѓ�����r�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h�d�    P��$V�`r3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    �m  j�D$ P�D$P���D$@�i���L$�D$4 �o  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�h�d�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     ��l  j �D$$P�D$P���D$D��h�����L$���D$8 �Pn  ��t:��r�t$@���   W��	���2�D$ P�F�D$<�����у��K��r�L$ ���   Q�@P���~ �t$D��rf��~@���   �D$$�	Pf�F�D$@�����у��ƋL$0d�    Y^[��0� �j�hd�    P��$V�`r3�P�D$,d�    ��r�t$<�D$     �D$(    ���   �L$ �@,Q�Ѓ��D$P�L$�D$8    �D$�  �D$    �D$    �k  j�D$ P�D$P���D$@�g���L$�D$4 �
m  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ��������j�hDd�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     ��j  j �D$$P�D$P���D$D��f�����L$���D$8 �@l  ��t3����r�L$ ���   Q�@8�Ѓ�����r�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�hod�    P��$V�`r3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    ��i  j�D$ P�D$P���D$@��e���L$�D$4 �Vk  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����j�h�d�    P��$SV�`r3�P�D$0d�    ���D$     �D$(    �D$P�L$�D$<    �D$�  �D$    �D$     �+i  j �D$$P�D$P���D$D�e�����L$���D$8 �j  ��t3����r�L$ ���   Q�@8�Ѓ�����r�D$ ���   P�	�D$<�����у��ƋL$0d�    Y^[��0�����������j�h�d�    P��$V�`r3�P�D$,d�    ��D$<�D$   �D$$�D$P�L$�D$8    �D$�  �D$    �D$    �<h  j�D$ P�D$P���D$@�4d���L$�D$4 �i  ��r�L$���   Q� �D$8�����Ѓ��L$,d�    Y^��0� ����������t��t��t3�ø   ���̡�rQ�@L�@L�Ѓ���������������̡�rQ�@L�@P�Ѓ���������������̡�r�t$�@L�t$�@TQ�Ѓ�� ���̡�r�t$�@LQ��  �Ѓ�� ����̡�r�t$�@LQ���   �Ѓ�� ����̡�rQ�@L�@X�Ѓ�����������������t$��r�t$�@L�t$�@\Q�Ѓ�� j�h�d�    P��0SVW�`r3�P�D$@d�    ��r�@L�@�Ћ؅�u�L$@d�    Y_^[��<� �L$�`���D$H    �D$(    �D$0    �D$4    �D$<    �D$8    �t$P�D$�D$0��r�\$(�@h]  �@0�L$�D$P�С�rj ���   j �@S���Ѕ���   ��rS�@L�@�Ћ�������   ����r���   �΋R(�ҋ��D$$Ph�   �t$0�  ����ts�L$<��tk��rj ���   ���   �ЋЅ�tP��rV���   �ʋ@<�С�r�L$<���   Q���   �Ѓ���t��rV�@@�@�Ѓ������`����+��rS�@@�@�С�r�L$@���   Q���   �Ѓ�3ۍL$$�D$H �e  �L$�D$H������^���ËL$@d�    Y_^[��<� ������������̡�rQ�@L�@`�Ѓ���������������̡�rQ�@L�@d�Ѓ���������������̡�r�t$�@LQ�@h�Ѓ�� �������̡�rQ�@L��D  �Ѓ������������̡�rQ�@L�@l�Ѓ���������������̡�r�t$�@LQ���   �Ѓ�� ����̡�r�@L�@����̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@L���   ��Y�������������̡�rQ�@L���   �Ѓ��������������t$��r�t$�@L�t$���   �t$�t$Q�Ѓ�� ������t$��r�t$�@L�t$���   Q�Ѓ�� ��������������t$��r�t$�@L�t$��   �t$Q�Ѓ�� ����������t$��r�t$�@L�t$��   Q�Ѓ�� ������������̡�r�@L��H  �࡜r�@L��L  �࡜r�@L��P  �࡜r�@L��T  �࡜r�@L��p  �࡜r�@L��t  �࡜r�@L���  �࡜r�@L���  �࡜r�@L���  �࡜r�@L���  ���T$ V�t$�D$hphPh@h0R�t$4�q�t$4�Q�t$4��r���@L�$�t$4���   VQ�Ѓ�4^�  ����̡�r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜rV�@�t$���   �6�Ѓ��    ^��������������̡�rV�@L�@�Ћ���u^á�rj �t$�@�t$��h  �t$V�Ѓ���u��rV�@@�@�Ѓ�3���^�������������̡�rj �H�t$�D$�� P�t$��h  �t$�Ѓ�������̡�r�@���   �࡜r�@L���   ���t$��r�t$�@�t$���   �t$ �t$ �t$ �t$�Ѓ��j�hd�    P�� V�`r3�P�D$(d�    �D$    �D$    �D$    �D$    �D$    �D$$    �D$     ��r�D$0    ���   ���   �ЉD$�t$8�D$0��t<��t8��rj�QLP���   ���ЋD$�D$ �D$Ph=���t$��	  ������   ��r�L$���   Q���   �D$4 �Ѓ��L$�D$    �D$0������  �ƋL$(d�    Y^��,������������j�hFd�    P�� V�`r3�P�D$(d�    �D$    �D$    �D$    �D$    �D$    �D$$    �D$     ��r�D$0    ���   ���   �ЉD$�t$8�D$0��t<��t8��rj�QLP���   ���ЋD$�D$ �D$Ph<���t$�  ������   ��r�L$���   Q���   �D$4 �Ѓ��L$�D$    �D$0�����   �ƋL$(d�    Y^��,�����������̡�r�@L���   �࡜r�@L���   �࡜r�@L��  �࡜r�@L��@  ���L$�� �������̋L$�t$��P��̋L$�t$��t$�P����������������t$�L$�t$��t$�t$�P������̡�r���   �AP���   ��Y�������̡�r�t$�@8Q�@D�Ѓ�� �������̡�r�@8�@<����̡�rV�@8�t$�@@�6�Ѓ��    ^���t$��r�t$�@8�t$�@�t$�t$�t$Q�Ѓ�� �����t$��r�t$�@8�t$�@�t$�t$Q�Ѓ�� �������̡�r�@8� �����̡�rV�@8�t$�@�6�Ѓ��    ^���t$��r�t$�@8�t$�@Q�Ѓ�� ��r�t$�@8�t$�@Q�Ѓ�� ���̡�rQ�@8�@�Ѓ���������������̡�r�t$�@8Q�@ �Ѓ�� ���������t$��r�t$�@8�t$�@$�t$�t$Q�Ѓ�� �������̡�r�t$�@8�t$�@(Q�Ѓ�� �����t$��r�t$�@8�t$�@,Q�Ѓ�� �t$��r�t$�@8�t$�@Q�Ѓ�� ��r�t$�@8�t$�@0Q�Ѓ�� �����t$��r�t$�@8�t$�@4Q�Ѓ�� ��r�t$�@8Q�@8�Ѓ�� �������̋L$��r�P�APP�A@P�A0P�A P�AP���   Q�t$�Ѓ����������������̡�r�@���   �࡜r�@���  �࡜r�@�@,����̡�r�@���  ��j�h�d�    PQV�`r3�P�D$d�    �D$    ��r�t$�@V�@�D$    �Ћ�rV�I�D$    �I8�D$   �у��ƋL$d�    Y^���������̡�r�@�@<����̡�r�@�@@����̡�r�@�@D����̡�r�@�@H����̡�r�@�@L����̡�r�@�@P����̡�r�@��<  �࡜r�@��,  ���t$��r�t$�@�t$���   �t$�t$h�2  �Ѓ����̡�r�@�@�����j�h�d�    P�� �`r3�P�D$$d�    ��r�L$�@Q�@�С�rj �@j��@�L$h@5Q���t$H�D$P�D$0P�D$L    ������r�L$$�@Q�@�D$P�С�r�L$8�@Q�@�С�r�L$<�@Q�@�D$X�����Ѓ�,�L$$d�    Y��,���������������̡�r�@���  �࡜r�@��8  ��j�h�d�    P��VW�`r3�P�D$ d�    �D$    ��r�L$�@Q��  �Ћ���r�|$4�IW�I�D$0   �ѡ�rW�@V�@�Ћ�r�D$ �IP�I�D$    �D$< �у��ǋL$ d�    Y_^�� ������������j�h(d�    P��VW�`r3�P�D$ d�    �D$    ��r�L$�@Q��  �Ћ���r�|$4�IW�I�D$0   �ѡ�rW�@V�@�Ћ�r�D$ �IP�I�D$    �D$< �у��ǋL$ d�    Y_^�� �����������̡�r�@��x  �࡜r�@��|  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@�@T����̡�r�@�@X����̡�r�@�@\����̡�r�@�@`����̡�r�@���  �࡜r�@�@d����̡�r�@�@h����̡�r�@�@l����̡�r�@�@p����̡�r�@�@t����̡�r�@��D  �࡜r�@��  �࡜r�@�@x����̡�r�@��@  ��j�hXd�    PQV�`r3�P�D$d�    �D$    �t$���D$    ��*����rV�I�t$$�I|�D$    �D$   �у��ƋL$d�    Y^������������̡�r�@���   �࡜r�@��d  �࡜r�@��h  �࡜r�@���  �࡜r�@���   ��j�h�d�    PQV�`r3�P�D$d�    �D$    �t$���D$    �sN����rV�I�D$    ���   �D$   �у��ƋL$d�    Y^�������������̡�r�@��`  �࡜r�@��  �࡜r���@�t$ ���   �L$Q�ЋL$$�~ f��~@f�A�~@f�A���� ��������������̡�r�@���  ���t$�D$��r���@�D$�D$���   �$�t$�Ѓ�����������̡�r�@���   �࡜r�@���   �࡜r�@���  �࡜r�@���  �࡜r�@��   �࡜r�@��  �࡜r�@��l  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@���  ��j�h�d�    P��VW�`r3�P�D$ d�    �t$4�D$    ��r�L$�@Q���  �Ћ���r�|$8�IW�I�D$4   �ѡ�rW�@V�@�Ћ�r�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� ��������j�h d�    P��VW�`r3�P�D$ d�    �t$4�D$    ��r�L$�@Q���  �Ћ���r�|$8�IW�I�D$4   �ѡ�rW�@V�@�Ћ�r�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� �������̡�r�@���  �࡜r�@���  ������r�T$�@R���   �T$R�T$RQ�����#D$���̃���r�T$�@R���   �T$R�T$RQ�����#D$���̃���r�$�@R���   �T$R�T$RQ�����#D$����̡�r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@���   �࡜r�@��  �࡜r�@��\  ��j�h8d�    P�� �`r3�P�D$$d�    �t$8�D$    ��r�L$�@Q��t  �Ѓ��t$4���D$0   ��'���L$�D$   �D$, � '���D$4�L$$d�    Y��,������������̡�r�@��H  �࡜r�@��T  �࡜r�@��p  �࡜r�@��8  ����  �`r3ĉ�$   ��$  P��$  �D$h   P�D0����x	=�  |'���rhH5�@hH  ��0  �Ѓ�Ƅ$�   ��r�$�@Q��4  hD5�Ћ�$  ��3���  ��  �������������������������t$$�D$�t$$�P�t$$��r�t$$�@0�t$$���   �t$$�t$$�t$$RQ�Ѓ�(�$ ��t$$�D$�t$$�P�t$$��r�t$$�@0�t$$���   �t$$�t$$�t$$RQ�Ѓ�(�$ ��t$$��r�t$$�@0�t$$���   �t$$�t$$�t$$�t$$�t$$�t$$Q�Ѓ�(�$ ����̡�rQ�@0���   �Ѓ������������̡�r�t$�@0�t$���   Q�Ѓ�� ��t$��r�t$�@0�t$���   �t$Q�Ѓ�� ��������̡�rQ�@0���   �Ѓ��������������t$��r�t$�@0�t$���   �t$Q�Ѓ�� ��������̡�r�@0���   �࡜rV�@0�t$���   �6�Ѓ��    ^���������������j�htd�    P��V�`r3�P�D$d�    �t$8�D$    ��r�t$8�@�t$8��X  �L$Q�ЋЋt$<j �    �F    ��rR���   V�@�D$@   �Ћ�r�D$(���   P�	�D$(   �D$D �у� �ƋL$d�    Y^�� ������������j�h�d�    P��(V�`r3�P�D$0d�    hLGOg�L$ �D$    ��E��j P�D$hicMCP�D$H   ��������L$�D$8�F����r�L$���   Q�@T�Ѓ���u�L$@�E���"��r�L$���   Q�@T�ЋL$D��P�E����r�D$���   P�	�D$   �D$< �ыD$D���L$0d�    Y^��4��������̡�r�@���  �࡜r�@���  �࡜r�@���  ��j�h�d�    P��VW�`r3�P�D$ d�    j �t$D�D$    �t$D��r�t$D�@�t$D��t  �L$$Q�Ћ���r�|$H�IW�I�D$D   �ѡ�rW�@V�@�Ћ�r�D$4�IP�I�D$4   �D$P �у�(�ǋL$ d�    Y_^�� ����������j�h0d�    P��V�`r3�P�D$d�    �t$<�D$    �t$<��r�t$<�@�t$<���  �L$Q�ЋЋt$@j �    �F    ��rR���   V�@�D$D   �Ћ�r�D$,���   P�	�D$,   �D$H �у�$�ƋL$d�    Y^�� ��������j�hSd�    P��$�`r3�P�D$(d�    ��r�@��p  �Ѕ���   h���L$�GC����r�t$8�@h���@4�L$�D$8    �С�r�t$<�@h���@4�L$��j �D$P�D$hicMCP������r�L$���   Q� �Ѓ��L$�D$0�����C���L$(d�    Y��0��������������j�h�d�    P��(VW�`r3�P�D$4d�    �D$    ��r�@��p  �Ѕ�u)��r�t$D�HV�I�у��ƋL$4d�    Y_^��4�h!���L$$�8B����r�t$H�@h!���@4�L$(�D$D   ��j �D$$P�D$hicMCP����P��r�D$P���   �@H�Ћ�r�|$X�IW�I���ы�rW�AV�@�Ћ�r�D$0���   P�	�D$0   �D$`�у�$�L$ �D$< ��A���ǋL$4d�    Y_^��4��������������j�h�d�    P��(VW�`r3�P�D$4d�    �D$    ��r�@��p  �Ѕ�u)��r�t$D�HV�I�у��ƋL$4d�    Y_^��4�h����L$$��@����r�t$H�@h����@4�L$(�D$D   ��j �D$$P�D$hicMCP�����P��r�D$P���   �@H�Ћ�r�|$X�IW�I���ы�rW�AV�@�Ћ�r�D$0���   P�	�D$0   �D$`�у�$�L$ �D$< �@���ǋL$4d�    Y_^��4��������������j�hd�    P��$V�`r3�P�D$,d�    ��r�@��p  �Ѕ�u�L$,d�    Y^��0�h#���L$��?����r�t$<�@h#���@4�L$ �D$<    ��j �D$P�D$hicMCP����P��r�D$H���   �@8�Ћ�r�����   �D$�	P�D$L �у��L$�D$4�����?���ƋL$,d�    Y^��0��������j�h1d�    P��$V�`r3�P�D$,d�    ��r�@��p  �Ѕ�u�L$,d�    Y^��0�hs���L$��>����r�t$<�@hs���@4�L$ �D$<    ��j �D$P�D$hicMCP�����P��r�D$H���   �@8�Ћ�r�����   �D$�	P�D$L �у��L$�D$4�����>���ƋL$,d�    Y^��0�������̡�r�@���  �࡜r�@���  �࡜r�@��@  ��V�t$���t��rQ�@��D  �Ѓ��    ^���������̡�r�@��H  �࡜r�@��L  �࡜r�@��P  �࡜r�@��T  �࡜r�@��X  �࡜r�@��\  �࡜r�@��d  �࡜r�@��h  �࡜r�@��l  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@��P  �࡜r�@���  ��j�hid�    P���`r3�P�D$d�    �t$0�D$    ��r�L$�@Q���  �Ѓ��L$,P�D$(   ��<���L$�D$   �D$$ ��<���D$,�L$d�    Y��$�������������̡�r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@���  �࡜r�@��l  �࡜r�@���  �࡜r�@���  �࡜r�@��$  �࡜r�@��(  �࡜r�@��,  �࡜r�@��0  �࡜r�@��<  �࡜r�@��  �࡜r�@��`  �࡜r�@��\  �࡜r�D$�@H���@�$Q�Ѓ�� �������������̡�rj �@HQ���   �Ѓ����������̡�r�t$�@Hj ���   Q�Ѓ�� ��̡�rj�@HQ���   �Ѓ����������̡�r�t$�@Hj���   Q�Ѓ�� ��̡�rj�@HQ���   �Ѓ���������̡�r�t$�@Hj���   Q�Ѓ�� ��̡�rQ�@H���  �Ѓ������������̡�r�t$�@HQ���  �Ѓ�� ����̡�r�t$�@HQ���  �Ѓ�� ����̡�r�t$�@HQ���  �Ѓ�� ����̡�r�t$�@H�t$��  Q�Ѓ�� ̡�r�t$�@H�t$��  Q�Ѓ�� ̡�rQ�@H���   �Ѓ�������������VW�t$��胐  ������t��r�t$�AHV���   W�Ѓ���_^� ���������VW�t$���t$���  ������t��r�t$�AHV���   W�Ѓ���_^� ����̡�r�t$�@H�t$���   Q�Ѓ�� ̡�r�t$�@H�t$���   Q�Ѓ�� ̡�r�t$�@HQ���   �Ѓ�� ����̡�rQ�@H���  �Ѓ��������������t$��r�t$�@H�t$���  �t$�t$Q�Ѓ�� �����j�h�d�    P��VW�`r3�P�D$ d�    ����rj �@Hh�  ���   W�Ѓ��|$0 ��   h�  �	�  ��������   ��rj �IHV���   W�у��L$��7����r�t$4�@h�  �@0�L$�D$0    �С�r�D$8�@���@,�$h�  �L$�С�rj �@@�L$�@(QV�Ѓ��L$�D$(�����7���   �L$ d�    Y_^�� � 3��L$ d�    Y_^�� � ������������̡�rQ�@H���   ��Y�������������̡�r�t$�@HQ���  �Ѓ�� ����̡�r�t$�@HQ���  �Ѓ�� ����̡�rQ�@H��4  �Ѓ������������̡�r�@H� �����̡�rV�@@�t$�@�6�Ѓ��    ^��S�\$U�l$V�}  W��u3��rS�@HW���   �Ѓ���u��rj�@HW���   �Ѓ���t�   �t$�E ����   ��rW�@H���   �Ѓ��|$( u!�t$$��rU�t$$�@HV���  SW�Ѓ��D��t@��I �t$$��rU�t$$�@HV���  SW�С�r�����   �΋@(�Ћ���uɋt$�}  u��rW�@H���   �Ѓ���t3���   �E ����rW�@Hu$���   �С�rS�@HW���   �Ѓ�_^][� ���   �С�r���|$( �@Hu!�t$$���  j �t$$VSW�Ѓ���_^][� � h  �Ћ����u_^][� ��r�΋��   �@x�Ћ�rP���   �͋B|�Ѕ�tP�t$$��rj �t$$�@HV���  SW�Ћȃ���t��rU���   �@H�С�r�΋��   �@(�Ћ���u�_^��][� ����t$��r�t$�@H�t$���  �t$�t$Q�Ѓ�� ����̡�rQ�@H���   ��Y�������������̡�rQ�@H���   �Ѓ������������̡�r�t$�@H�t$���   Q�Ѓ�� ̡�rQ�@H���   ��Y�������������̡�rQ�@H��t  ��Y�������������̡�rQ�@H��P  �Ѓ������������̡�rQ�@H��T  �Ѓ������������̡�rQ�@H��X  �Ѓ������������̡�r���@HQ��\  �L$Q�ЋL$$�~ f��~@f�A�~@f�A���� � ��������������̡�rQ�@H��`  �Ѓ������������̡�r�t$�@HQ��d  �Ѓ�� ����̡�r�D$�@H����h  �$Q�Ѓ�� ����������̡�r�D$�@H����t  �$Q�Ѓ�� ����������̡�r�D$�@H����l  �$Q�Ѓ�� ����������̡�r�t$�@HQ��p  �Ѓ�� ������t$��r�t$�@H�t$���  �t$Q�Ѓ�� ����������t$��r�t$�@H�t$���  �t$�t$�t$Q�Ѓ�� ̡�rh�  �@H� �Ѓ������������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@H���   �Ѓ������������̡�rQ�@H���   �Ѓ������������̡�r�t$�@HQ���   �Ѓ�� ����̡�r�t$�@HQ���   �Ѓ�� ����̡�r�t$�@H�t$��   Q�Ѓ�� ��t$��r�D$�@H�����  �$Q�Ѓ�� ������̡�rV�@Hh  � �Ћ�������   �t$h�  �#�  �Ѓ���t^��rj �AHR���   V���t$h(  ���  �Ѓ���t2��rj �AHR���   V�С�r�����   j �@j���Ћ�^á�rV�@@�@�Ѓ�3�^�������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@H��  �Ѓ������������̡�rQ�@H��  �Ѓ������������̡�rQ�@H���  �Ѓ������������̡�rQ�@H���  �Ѓ������������̡�rQ�@H���  �Ѓ������������̡�r�t$�@H�t$��  Q�Ѓ�� ��t$��r�t$�@H�t$��   Q�Ѓ�� ��������������t$��r�t$�@H�t$��|  �t$Q�Ѓ�� ��������̋D$V���u��r�@H���  �'��u��r�@H���  ���u(��r�@H���  V�Ѓ���tP�t$���   ^� 3�^� ������������̃�SVW���ӏ  �؅���   �|$$����   ��rj �AHh�  ��p  V�Ѓ��D$��u_^��[��� U3�ωl$�`�  ����   ���    �D$P�D$PU����  ��tf�t$;t$\�l$������u����ɋD�;D�t.��r�Hl����P�D$(�p�A�ЋD������tP����  F;t$~��l$�|$(E�ωl$�ȋ  ;��p���]_^��[��� _^3�[��� ��������̃���rU�@Hj ��p  ��h�  U�l$�Ѓ��D$��u]��� �D$W��u��r�@H���  �+��u��r�@H���  ����Z  ��r�@H���  U�Ћ������<  S��菋  ��rh�  �@H3ۋ��   U�\$(�Ѓ�����   �l$V�s����r�L$�@lS�q�@�Ћ؃�����   ��r�s�I\�t$$�I,�у���t�F�P��贊  ��r�s�@\�t$$�@,�Ѓ���t�F�P��莊  �E ;Et#��r�s�@\�t$$�@,�Ѓ���tV���c�  ��r�s�@\�t$$�@,�Ѓ���t�FP���=�  ��r�\$$�@Hh�  �t$���   C�\$,�����Ѓ�;�����^[_�   ]��� _3�]��� ̡�rQ�@H���  �Ѓ������������̡�r�t$�@H�t$���  Q�Ѓ�� ��t$��r�t$�@H�t$���  Q�Ѓ�� ������������̡�rQ�@H���  �Ѓ������������̡�rQ�@H���  �Ѓ������������̡�r�t$�@HQ��  �Ѓ�� ����̡�r�t$�@HQ��  �Ѓ�� ����̡�rQ�@H��  �Ѓ������������̡�r�t$�@HQ��  �Ѓ�� ����̡�rQ�@H��T  �Ѓ������������̡�r�t$�@H�t$��  Q�Ѓ�� ̡�r�t$�@HQ��8  �Ѓ�� ����̡�r�t$�@HQ��<  �Ѓ�� ������t$��r�t$�@H�t$��@  Q�Ѓ�� ������������̡�r�t$�@HQ���  �Ѓ�� ����̡�r�t$�@HQ��H  �Ѓ�� ����̡�rQ�@H��L  ��Y�������������̡�rV�@Hh�  � �Ћ�����u^á�r�t$�@H�t$��  V�Ѓ���u��rV�@@�@�Ѓ�3���^������������̡�rV�@@�t$�@�6�Ѓ��    ^���t$��r�t$�@H�t$��   Q�Ѓ�� ������������̡�r�D$�@H����$  �$Q�Ѓ�� ����������̡�rQ�@H��(  �Ѓ������������̡�r�t$�@H�t$��,  Q�Ѓ�� ̡�r�@H��  �࡜r�@H��  �࡜rV�@@��@,WV�Ћ�r���ȋBj ���   h�  �Ћ�rh�  �IHV���   ���у���
��t_3�^Ë�_^�̡�rQ�@@�@,�Ћ�r���ЋAj ���   h�  ������̡�r�D$�@H����  �t$,�t$,���$Q�L$Q�ЋL$4�~ f��~@f�A�~@f�A����0� ��������̡�r�D$�@H����  �t$,�t$,���$Q�L$Q�ЋL$4�~ f��~@f�A�~@f�A����0� ��������̡�rQ�@H���  �Ѓ������������̡�r�t$�@H�t$��8  Q�Ѓ�� ��t$��r�D$�@H����0  �$�t$Q�Ѓ�� ��̡�r�@H�@����̡�rV�@@�t$�@�6�Ѓ��    ^���t$�D$�t$��r���@H�$�t$���   �t$�t$�Ѓ�������������t$�D$��r���@H�$�t$���   �t$�t$�Ѓ�����������������    ���������̡�rj�@H�1��|  �Ѓ���������̡�rV�@H�t$��x  ����3Ƀ������^��� ������̡�rj �@H�1��|  �Ѓ����������fnD$�L$����YD$�Xh6�,�;�}���;D$OD$���������������̃�D��rS�@HV���   W�|$Th�  W�Ћ�r3��IHV���   ��h�  W�\$H�у��D$H�t$�t$�t$��u
_^�C[��Dá�rU���   �ϋ@��=�  ��r�@  �@Hj ���   h:  W�Ћ�rh�  �IHW���   �D$0�ы�r3�IHU���   h�  W�D$H�ы�r�؋IHW��  �\$D�ы�rW�IH�D$d���  �у�(3��D$@�D$Pd69t$(�|   �K�ً��D$<��tPj�W��讣  ���tA�L$@�@�|� ���L$H~�� ��%�������;�u&�*�  �L$H;�O���  ���;Cu�����G��;|$(|��\$ �D$�|$X���|   j W����  ����  �L$�  ��t]�L$�z  �L$8;�uL��r�I�@h�5���  ��h�  Q�L$T�Ѓ��D$����  �L$P�t$LP�H  P�  ���D$8h�5�@��r���@h�  ���  Q�L$T�Ѓ��D$���@  �T$L��t�L$H��tQRP��  ����~-��rh�5�@h�  ���   ��U�Ѓ��D$����  ��rj��@HV��  W�Ѓ�����  �l$��t!jW����~  ����  ���~  ���D$,�3��t$,��rj �@Hh�  ���   W�Ћ�3�3���T$�l$$�D$49D$(�h  �{�|$8�L$<���u  j�P蛡  ����`  �L$@�@�|� �4��t$H~�� ��%�������9D$4��  ���۝  3�3��D$L�D$0    9^��   �l$ ��������Шtm�D$������������������D$���T��N�D$�L��D$�J�L��N�D$�L���D$�J�L��N�D$�t$H�L���D$�J�L��C;^�y����l$$���7  �Ǚ+�j��P�t$�L$\�T�  �\$�L$,�m    �3��Ë�+ÉD$D�T$H��;D$L�  �D$����t3�D$�l$D�[�~�f�*�~D�f�D*�~D��ŋl$$f�D�D$�[�~�f��~D�f�B�~D�f�B;�}_�D$9�uR�L�����������w4�$�E�L$ ��,��"�L$ ��l���L$ ��l��
�L$ ��l���;�|��T$H�D$0�L$,E��@�l$$�T$H�D$0;�����;D$L�-  �|$8�T$�D$4�t$,@���D$4�|$8;D$(������D$P�4����D$P�*������  �T$��L$3�;G�Å���   �m    ōƋG��@�~�f��~D�f�B�~D�f�B�G��@�D$�~�f�B�~D�f�B �~D�f�B(��T$�@�D$�~ȍȍm    �f�D�0�~Af�D�8�~Af�D�@��t7�G�@�D$�~ȍȍm    �f�D�H�~Af�D�P�~Af�D�X�G��@�D$�~ȍȍm    �f���~Af�D��~Af�D��G��o��@�D$E�~ȍȍm    �f���~Af�D��~Af�D���o��@�D$E�~ȍȍm    �f���~Af�D��~Af�D��/E�l$$��tC�G�@�D$�~ȍȍm    �f���~Af�D��~Af�D��oE�l$$�������G������D$P�-����D$P�#����D$P������3�]_^[��DË��   �ϋ@��=  ��  ��rj �@Hh(  ���   W�Ћ�rh(  �IHW���   ���ы��3ɉl$D��~�d$ �˅�t�|� �4Vu���A;�|�D$8h6�@��r���@hK  ���  Q�L$\�Ћȃ��L$����   �T$L��t�D$P��tPRQ���  ����rh,6�@��    ���  hP  Q�Ћȃ��L$$��tW��t��    ��tPSQ趷  ����r�ƋIH���   +���PVW�D$L�у���u!�D$P������D$(P������]_^3�[��Dá�rj �@Hh�  ���   W�Ћ�rj �IHh(  ���   W�D$d��3�3ۃ���3҉L$P�t$H�\$8���#  �|$$���$    ��߅���   3��~y�L$L�R�4v�]�����D$C�~f��~Df�A�~Df�A�D$���~Df�A�~D f�A �~D(�D$8f�A(�|$$E�I0�v;�|��t$H�؃|� tg�|$L�.�@�D$�~ȍȍRBf���~Af�D��~Af�D��D$�v�~ȍȍRBf���~Af�D��~Af�D��|$$4ߋl$D�t$HC�\$8;�������L$P�T$@3���~��D�    ��   @;�|�D$$P�������D$P�������   ]_^[��DÐI?T?`?l?�����t$�D$��r���@H�$�t$���  �t$�Ѓ���̡�r�@H���  �࡜r�@H���  ���t$,�D$(��r���@H�$�t$,���  �t$,�t$,�t$,�t$,�t$,�t$,�t$,�Ѓ�,����������̡�r�@H���  �࡜r�@H���  ���t$,�D$�t$,��r�t$,�@H�t$,��P  �t$,���D$�D$0�$�t$,�t$,�Ѓ�,��������X6�A    ����q�X6��r�@l�@��Y��������̡�rV�@l��@�v�ЋL$����u	�   ^� �t$��r�t$�@lQ�t$� ��3Ƀ������F^��� ������������̋I��u3�á�rQ�@l�@�Ѓ�����̃���r�$�@lR�@�T$R�t$�t$�q�ЋL$�T$(��;�u	�$��� ���9$D���� ����̡�r�@H���   �࡜r�@H���  ������r�L$�@�����   W��$�t$���$�D$�$f/�w�D$f/�w(���r�L$�@���@,�$�t$�Ѓ�������̃�0��rW��$Q�t$<�D$�D$�D$�@�L$ ���   Q�L$@���~X�D$<f/��~ �~P�L$Dv(��	f/�v(�f/�v(��	f/�v(�f/�wf/�v(��(ġ�r�$�T$�\$�@�$�@HQ�t$<�L$<�Ѓ�0���̡�r�@H��0  ���������������������������������̡�r�@H���  �࡜r�@H���  ���t$,��r�t$,�@H�t$,���  �t$,�t$,�t$,�t$,�t$,�t$,�t$,�t$,Q�Ѓ�0�, ��������������t$,��r�t$,�@H�t$,���  �t$,�t$,�t$,�t$,�t$,�t$,�t$,�t$,Q�Ѓ�0�, ������������̡�rQ�@H��,  �Ѓ������������̡�r�t$�@HQ��X  �Ѓ�� ����̡�rQ�@H��\  �Ѓ������������̡�rQ�@H�t$���   �t$�Ѓ�� ̋D$��t�L$��t�T$��tRPQ誰  ���������������V���v�X6��r�@l�@�Ѓ��D$t	V�g�������^� �������������̋D$�L$� +� ̸   � ��������3�� �����������3�� ����������̸   @� ��������3�� ����������̸   � ��������Q��r�t$�H�D$    �I�ыD$��� �����������̸   � �������́��   V��$�   ��u
3�^���   �h�   �D$j P�k�  ��$�   �D$P��$�   �D$T��$�   h�   �D$�D$P��$�   �t$<��$�   �D$$�8 j�D$lk �D$piO�D$tnOǄ$�   'k �D$|"k Ǆ$�   k Ǆ$�   dOǄ$�   sO蛿���� ^���   Á��   h�   �D$j P豮  ��$�   h�   �D$P�D$P��$�   �D$8    ��$�   j�G������   �j�h�d�    P��   SVW�`r3�P��$�   d�    3ۉ\$��$�   3���$�   ����  ��r��$�   �@�@<�Ѕ��B  �u3  �D$Ƅ$�   ���  ��$�   P�L$L�p�����r�L$�@Q�@Ƅ$�   �D$   �С�rV�@j��@�L$(hp6Q�Ѓ��D$P�L$0Ǆ$�      �D$   ������$�   PǄ$�      �D$   ����L$0QP��$�   PǄ$�      �D$    ������L$XQP�D$|PǄ$�      �D$,   �������L$Vj��?   PǄ$�      �\$�/  �D$��t�D$ Ǆ$�      �� t��ߍL$d�\$�T���Ǆ$�      ��t��$�   �\$�1���Ǆ$�      ��t�����$�   �\$����Ǆ$�      ��t����L$,�\$�����Ǆ$�      ��t��r�L$�@����@Q�\$�Ѓ�Ǆ$�      ��t	�L$H�����|$ t+W��$�   �t$ ��$�   ��$�   ��$�   �\��������D$PƄ$�    �U1  ���D$    �)W��$�   j ��$�   ��$�   ��$�   ����������r��$�   �IP�IǄ$�   �����у��Ƌ�$�   d�    Y_^[�Ĵ   �V��V��0  ���    ^Ë�`��`��`��`���������    �A    �A    �A    �����V��~ u=���t��rQ�@<�@�Ѓ��    W�~��t���k���W��������F    _^���������j�h�d�    P��V�`r3�P�D$$d�    ��D$P�@����P���D$0    �-   �L$���D$,����������ƋL$$d�    Y^��(��������j�h�d�    PQV�`r3�P�D$d�    ��~ uWht6j;h�rj��������D$�D$    ��t�t$�������3��D$�����F��u�L$d�    Y^��� �~ t3�9�"��r�t$�@<� �Ћȃ�3���F   �����L$d�    Y^��� �����������V���F   ��r�@<�@��3Ʌ����^��������������̋	��r��u�@� � �@<�t$�@Q�Ѓ�� ���������̃y t�   ËQ��u3�á�rR�@<�1�@�Ѓ��������V��~ u=���t��rQ�@<�@�Ѓ��    W�~��t���K���W��������F    _^��������̋|r��r��u�@� Ë@<�t$�@Q�Ѓ������������j�h@d�    P��(SV�`r3�P�D$4d�    �D$    �|r��u��r�A�0���r�t$H�@<Q�@�Ћ�r�����I�D$�IP�ѡ�r�L$�@Q�@V�С�r�L$0�@Q�@�D$L   �С�rj �@j��@�L$<h�6Q�Ѓ� ��rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@��tA�t$D�@V�Ћ�r�D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С�rj��@j��t$T�@L�t$�L$$�С�r�t$D�@V�@�С�r�L$�@V�@Q�Ћ�r�D$ �IP�I�D$    �D$L �у��ƋL$4d�    Y^[��4��j�h�d�    P��(SV�`r3�P�D$4d�    �D$    �|r��u��r�A�0���r�t$H�@<Q�@�Ћ�r�����I�D$�IP�ѡ�r�L$�@Q�@V�С�r�L$0�@Q�@�D$L   �С�rj �@j��@�L$<h�6Q�Ѓ� ��rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@��tA�t$D�@V�Ћ�r�D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С�rj��@j��t$T�@L�t$�L$$�С�r�L$$�@Q�@�С�rj �@j��@�L$0h�6Q�Ѓ���rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@��t�t$D�@V�������@Hj�t$�L$�С�rj��@j��t$X�@L�t$�L$$�С�r�t$D�@V�@�С�r�L$�@V�@Q�Ћ�r�D$ �IP�I�D$    �D$L �у��ƋL$4d�    Y^[��4����������j�h�d�    P��(SV�`r3�P�D$4d�    �D$    �|r��u��r�A�0���r�t$H�@<Q�@�Ћ�r�����I�D$�IP�ѡ�r�L$�@Q�@V�С�r�L$0�@Q�@�D$L   �С�rj �@j��@�L$<h�6Q�Ѓ� ��rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@��tA�t$D�@V�Ћ�r�D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С�rj��@j��t$T�@L�t$�L$$�С�r�L$$�@Q�@�С�rj �@j��@�L$0h�6Q�Ѓ���rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@��t�t$D�@V�������@Hj�t$�L$�С�rj��@j��t$X�@L�t$�L$$�С�r�L$$�@Q�@�С�rj �@j��@�L$0h�6Q�Ѓ���rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@���D����@Hj�t$�L$�С�rj��@j��t$\�@L�t$�L$$�С�r�t$D�@V�@�С�r�L$�@V�@Q�Ћ�r�D$ �IP�I�D$    �\$L�у��ƋL$4d�    Y^[��4��������������j�h<d�    P��(SV�`r3�P�D$4d�    �D$    �|r��u��r�A�0���r�t$H�@<Q�@�Ћ�r�����I�D$�IP�ѡ�r�L$�@Q�@V�С�r�L$0�@Q�@�D$L   �С�rj �@j��@�L$<h�6Q�Ѓ� ��rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@��tA�t$D�@V�Ћ�r�D$�IP�I�D$   �D$D �у��ƋL$4d�    Y^[��4Ë@Hj�t$�L$�С�rj��@j��t$T�@L�t$�L$$�С�r�L$$�@Q�@�С�rj �@j��@�L$0h�6Q�Ѓ���rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@��t�t$D�@V�������@Hj�t$�L$�С�rj��@j��t$X�@L�t$�L$$�С�r�L$$�@Q�@�С�rj �@j��@�L$0h�6Q�Ѓ���rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@���D����@Hj�t$�L$�С�rj��@j��t$\�@L�t$�L$$�С�r�L$$�@Q�@�С�rj �@j��@�L$0h�6Q�Ѓ���rj �@�L$�@@Q�L$,Q�L$ �D$H�Ѕ���r�L$$�@Q�@���D$@�С�r���@��������@Hj�t$�L$�С�rj��@j��t$`�@L�t$�L$$�С�r�t$D�@V�@�С�r�L$�@V�@Q�Ћ�r�D$ �IP�I�D$    �\$L�у��ƋL$4d�    Y^[��4ËD$�|r��EȉL$��  �������̡�r�@<�@����̋D$����u���VP�L$�S  �D$P�D$P�L$�D$    �D$    �S  ����   �t$��$    �D$��tB��t=��uZ��r�t$���   �@H�Ћ�r�ЋA���@xV���Ѕ�u,�   ^��á�r�t$���   �@T��VP�J�������uԍD$P�D$P�L$� S  ���x���3�^����j�h�d�    P��HSUVW�`r3�P�D$\d�    3ۉ\$��r�L$,�@Q�@�С�rS�@j��@�L$8h�6Q�С�r�L$@�@<Q�@�\$|�Ћ�r���I�D$D�IPǄ$�   �����у���u3��L$\d�    Y_^][��T�V�L$(3��R  �D$P�D$$P�L$,�ER  ���  �l$l���$    �|$ ��   ��r�t$���   �@T�Ћ�����tc��r�D$<�IP�I�у��D$<Pj�D$T��P���D$p   �\$$� ~���Ћ�r���AU�@x���D$h   �\$���D$��t�D$ �D$d   ��t��r�L$L�@����@Q�\$�Ѓ��D$d������t��r�L$<�@Q�@����Ѓ��|$ u�D$P�D$$P�L$,�8Q  ��� �����|$�ǋL$\d�    Y_^][��T�����j�h�d�    P��DSUVW�`r3�P�D$Xd�    �t$l3ۉ\$��u|��r�L$(�@Q�@�С�rV�@j��@�L$4h�6Q�С�r�L$<�@<Q�@�t$x�Ћ�r���I�D$@�IP�D$|�����у���u3��L$Xd�    Y_^][��P�V�L$$3��P  �D$P�D$ P�L$(�@P  ����   �|$h�d$ �D$����   ��r�t$���   �@T�Ћ�����tc��r�D$8�IP�I�у��D$8Pj�D$P��P���D$l   �\$$��{���Ћ�r���AW�@x���D$d   �\$���D$l��t�D$l �D$`   ��t��r�L$H�@����@Q�\$�Ѓ��D$`������t��r�L$8�@Q�@����Ѓ��|$l tR�l$�ŋL$Xd�    Y_^][��PÃ�u3�L$��t+��rQ���   �@H�Ћ�r�ЋA���@xW���Ѕ�t��D$P�D$ P�L$(��N  �����������������̡�r�@<�@����̃=�r uK�|r��t��rQ�@<�@�Ѓ��|r    V�5�r��t�������V�Z�������r    ^�����������̋D$V�0W�9;�t_3�^� �P��u��u9pu9qu��u�9yu�_�B^� S�Y��u!��u9yu��u2��u.9pu)[_�   ^� ��t��t;�u�P��t�A��t�;�t�[_3�^� �������t$�g������@� ���������������Vh�rj\hD ��輂  ����t�@\��tV�Ѓ���^�����Vh�rj\hD ��茂  ����t3�@\��t,V��h�rjxhD �j�  ����t�@x��t
V�t$�Ѓ���^� �����������̃�Vh�rj\hD ���)�  ����tL�@\��tEV�ЋD$h�rjdhD �D$�D$    �D$    ��  ����t�@d��t�L$QV�Ѓ���^��� �������������Vh�rj\hD ��謁  ����t3�@\��t,V��h�rjdhD 芁  ����t�@d��t
�t$V�Ѓ���^� ������������Vh�rj\hD ���L�  ����t\�@\��tUV��h�rjdhD �*�  ����t�@d��t
�t$V�Ѓ�h�rjhhD ��  ����t�@h��t
�t$V�Ѓ���^� ���Vh�rj\hD ���̀  ������   �@\��t~V��h�rjdhD 覀  ����t�@d��t
�t$V�Ѓ�h�rjhhD �}�  ����t�@h��t
�t$V�Ѓ�h�rjhhD �T�  ����t�@h��t
�t$V�Ѓ���^� ������Vh�rj`hD ����  ����t�@`��tV�Ѓ�^�������Vh�rjdhD ����  ����t�@d��t
�t$V�Ѓ�^� Vh�rjhhD ���  ����t�@h��t
�t$V�Ѓ�^� Vh�rjlhD ���  ����t�@l��tV�Ѓ�^�������Vh�rjphD ���\  ����t�@p��t�t$V�Ѓ�^� ��r^� �������Vh�rjxhD ���  ����t�@x��t
V�t$�Ѓ���^� ��������������Vh�rj|hD ����~  ����t�@|��tV�t$�Ѓ�^� 3�^� ����������Vh�rj|hD ���~  ����t�@|��tV�t$�Ѓ����@^� �   ^� ��j�h1d�    P��V�`r3�P�D$d�    ��h�rjthD �D$    �1~  ����tu�@t��tn�t$(�L$VQ�Ѓ��t$$P���D$    �`���h�rj`hD �D$   �D$( ��}  ����tv�H`��to�D$P�у��ƋL$d�    Y^��� h�rj\hD �}  �t$0����t4�@\��t-V��h�rjdhD �~}  ����t�@d��th�rV�Ѓ��ƋL$d�    Y^��� Vh�rh�   hD ���9}  ����t���   ��t�t$V�Ѓ�^� 3�^� ����Vh�rh�   hD ����|  ����t���   ��t�t$V�Ѓ�^� 3�^� ����VW��3����$    �h�rjphD �|  ����t�@p��t	VW�Ѓ����r�8 tF��_��^�������SU�l$V��3�W�d$ h�rjphD �_|  ����t�@p��t	VS�Ѓ����r�8 tnh�rjphD �-|  ����t�@p��tVU�Ѓ������rh�rjphD ��{  ����t�@p��t	VS�Ѓ����rW���Z�����tF�`����D$_��t�0��~=h�rjphD �{  ����t�@p��t	VS�Ѓ����r�8 u^]�   [� ^]3�[� �����������̃�Vh�rh�   hD ���V{  ����t?���   ��t5�t$�L$VQ��h�rj`hD �({  ����t�@`��t
�L$Q�Ѓ���^��� �������j�hmd�    P��V�`r3�P�D$d�    h�rh�   hD �D$    ��z  ����ty���   ��to�t$,�L$�t$,Q�Ѓ��t$$P���D$    �����h�rj`hD �D$   �D$( �kz  ����ts�H`��tl�D$P�у��ƋL$d�    Y^���h�rj\hD �/z  �t$0����t3�@\��t,V��h�rjxhD �	z  ����t�@x��t
V�t$,�Ѓ��ƋL$d�    Y^����������������̋���������������h�rjhD �y  ����t	�@��t��3��������������V�t$�> t+h�rjhD �uy  ����t�@��tV�Ѓ��    ^���������̃|$ W��t1h�rjhD �5y  ����t�@��t�t$�t$W�Ѓ�_� 3�_� ���������������Vh�rjhD ����x  ����t�@��t�t$V�Ѓ�^� 3�^� ����������Vh�rjhD ���x  ����t�@��t�t$V�Ѓ�^� 3�^� ����������Vh�rj hD ���lx  ����t�@ ��tV�Ѓ�^�3�^���Vh�rj$hD ���<x  ����t�@$��tV�Ѓ�^�3�^���Vh�rj(hD ���x  ����t�@(��t�t$�t$�t$V�Ѓ�^� 3�^� ��Vh�rj,hD ����w  ����t�@,��t�t$�t$V�Ѓ�^� 3�^� ������Vh�rj(hD ���w  ����t�@0��t�t$�t$�t$V�Ѓ�^� 3�^� ��Vh�rj4hD ���Lw  ����t�@4��tV�Ѓ�^�3�^���Vh�rj8hD ���w  ����t!�@8��t�t$�t$�t$�t$V�Ѓ�^� 3�^� ��������������Vh�rj<hD ����v  ����t�@<��t
�t$V�Ѓ�^� Vh�rh�   hD ���v  ����u^� �t$���   V�Ѓ�^� ����������Vh�rh�   hD ���Yv  ����u^� �t$���   V�Ѓ�^� ����������Vh�rh�   hD ���v  ����u^� �t$���   V�Ѓ�^� ����������Vh�rh�   hD ����u  ����t�t$���   �t$�t$V�Ѓ�^� ������Vh�rjDhD ���u  ����t�@D��tV�Ѓ�^�3�^���Vh�rjHhD ���lu  ����t�t$�@HV�Ѓ�^� ����Vh�rjLhD ���<u  ����u^� �t$�@LV�Ѓ�^� Vh�rjPhD ���u  ����u^� �t$�@P�t$V�Ѓ�^� ������������Vh�rh�   hD ����t  ����u^� �t$���   �t$�t$V�Ѓ�^� ��Vh�rh�   hD ���t  ����u^� �t$���   �t$�t$�t$�t$V�Ѓ�^� ����������Vh�rjThD ���<t  ����u^Ë@TV�Ѓ�^���������Vh�rjXhD ���t  ����t�t$�@XV�Ѓ�^� ����j�h�d�    P��V�`r3�P�D$ d�    ��h�rh�   hD �D$    �s  ����t~���   ��tt�t$4�L$Q���Ћt$0P���D$,   �����h�rj`hD �D$   �D$4 �^s  ������   �H`����   �D$P�у��ƋL$ d�    Y^��$� h�rj\hD �D$     �D$$    �D$(    � s  �t$<����t4�@\��t-V��h�rjdhD ��r  ����t�@d��t�L$QV�Ѓ��ƋL$ d�    Y^��$� ������������Vh�rh�   hD ���r  ����t���   ��t�t$���t$�t$��^� 3�^� ��������������Vh�rh�   hD ���9r  ����t���   ��t�t$����^� 3�^� ������Vh�rh�   hD ����q  ����t���   ��t�t$����^� 3�^� ������Vh�rh�   hD ���q  ����t���   ��t�t$����^� 3�^� ������Vh�rh�   hD ���yq  ����t���   ��t��^��3�^����������������Vh�rh�   hD ���9q  ����t���   ��t�t$���t$�t$��^� 3�^� ��������������Vh�rh�   hD ����p  ����t���   ��t�t$����^� ������������Vh�rh�   hD ���p  ����t���   ��t�t$���t$�t$��^� 3�^� ��������������Vh�rh�   hD ���Yp  ����t���   ��t��^��3�^����������������h�rjhD �p  ����t	�@��t��3��������������j�h�d�    P��VW�`r3�P�D$ d�    h�rh�   hD �D$    �o  ����u)��r�t$0�HV�I�у��ƋL$ d�    Y_^�� ��t$4���   �L$Q�Ћ���r�|$8�IW�I�D$4   �ѡ�rW�@V�@�Ћ�r�D$$�IP�I�D$$   �D$@ �у��ǋL$ d�    Y_^�� ������������h�r�t$hD ��n  �����������̋D$��r� ����̡�r�@��   �࡜rV�@�t$��$  �6�Ѓ��    ^��������������̡�rV�@��(  V�t$�Ѓ���^� ��������������̡�rQ�@�t$��,  �Ѓ�� ����̡�rQ�@�t$��,  �Ѓ����@� �D$��t�P�3ҡ�rR�@Q��8  �Ѓ�� ��������̡�r�t$�@Q��<  �Ѓ�� ������t$��r�t$�@�t$��@  Q�Ѓ�� ������������̡�r�t$�@�t$��D  Q�Ѓ�� ̡�r�t$�@Q��H  �Ѓ�� �����j�h!d�    P��VW�`r3�P�D$ d�    �t$4�D$    ��rQ�@�L$��L  Q�Ћ���r�|$<�IW�I�D$8   �ѡ�rW�@V�@�Ћ�r�D$(�IP�I�D$(   �D$D �у��ǋL$ d�    Y_^�� � ���̡�rQ�@��T  �Ѓ������������̡�rQ�@��P  �Ѓ������������̡�r�t$�@Q��X  �Ѓ�� ����̡�r�t$�@Q��l  �Ѓ�� ����̡�r�@��0  �࡜r�@��4  �࡜r�@��p  �࡜r�@��t  �࡜r�@��\  �࡜rV�@�t$��`  �6�Ѓ��    ^����������������t$��r�t$�@�t$��d  �t$�t$Q�Ѓ�� ������t$��r�t$�@�t$��h  �t$�t$Q�Ѓ�� ����̡�rQ�@�@�Ѓ�����������������t$��r�t$�@�t$�@X�t$Q�Ѓ�� �����������̡�r�t$�@Q�@\�Ѓ�� �������̡�rQ�@�@ ��Y�j�hDd�    P��V�`r3�P�D$d�    ��rh�  �@Q���   �L$Q��P��r�D$0    ���   �@8�Ћ�r�����   �D$�	P�D$4�����у��ƋL$d�    Y^����̡�r�@��   ���t$��r�t$�@�t$�@Q�Ѓ�� �t$��r�t$�@�t$���   �t$Q�Ѓ�� ��������̡�r�@�@$������t$��r�t$�@�t$�@(�t$Q�Ѓ�� �������������t$��r�t$�@�t$�@,�t$Q�Ѓ�� �������������t$$��r�t$$�@�t$$�@`�t$$�t$$�t$$�t$$�t$$�t$$Q�Ѓ�(�$ �������̡�rV�@W�@��W�Ћ�rW�J���I���t$��r�t$�Q�t$�N�QHP�B4j j W�Ѓ�(_^� �t$��r�t$�@�t$�@4�t$�t$�t$�t$Q�Ѓ� � ��r�t$�@�t$�@@Q�Ѓ�� ���̡�r�t$�@Q�@D�Ѓ�� �������̡�rQ�@�@L�Ѓ���������������̡�rQ�@�@L�Ѓ���������������̡�rQ�@�@P�Ѓ���������������̡�r�t$�@Q�@T�Ѓ�� �������̡�r�t$�@Q�@T�Ѓ�� �������̡�rQ�@�@h�Ѓ���������������̡�r�t$�@�t$���   Q�Ѓ�� �j�h�d�    P��V�`r3�P�D$d�    �t$4�D$    ��r�t$4�@Q���   �L$Q�ЋЋt$<j �    �F    ��rR���   V�@�D$@   �Ћ�r�D$(���   P�	�D$(   �D$D �у� �ƋL$d�    Y^�� � �����������̡�r�@� �����̡�rV�@�t$�@�6�Ѓ��    ^���t$��r�t$�@�t$���   �t$�t$Q�Ѓ�� ����̡�rV�@�t$�@�6�Ѓ��    ^��QVW�|$����m  ��rV�@�@h�Ѓ�����ru �@h|7��0  h�  �Ѓ�_3�^Y� �L$Q�L$Q�t$�D$    �@V���   �Ѓ���tϋL$3���~�I �D$����tP���k  �L$F;�|�D$P�ʳ�����   _^Y� ������������QVW�|$�����l  ��rV�@�@h�Ѓ�����ru �@h�7��0  h�  �Ѓ�_3�^Y� �L$Q�L$Q�t$�D$    �@V���   �Ѓ���tσ|$ t�3�9t$~5�D$����t#��rQ�@�@h�Ѓ���t�D$���4��j  F;t$|ˍD$P�������   _^Y� ̡�r�@��x  �࡜r�@��|  �࡜rQ�@���   �Ѓ������������̡�r�t$�@Q���   �Ѓ�� ����̡�r�@���   �࡜rV�@�t$���   �6�Ѓ��    ^���������������VW���O�t���W�f�G f�G(f�G0f�G8f�G@f�GHf�GPf�GX�    �G`    �Gd    �Gh    �Gp�Gx�����G|   ��_^�������j�h�d�    PQV�`r3�P�D$d�    ��t$�D$    �k   �N�D$����軸���L$d�    Y^�������������W��    �A`    �Ad    �Ah    �Ap�Ax�����A|   ���������������SW�����t7��迴���xP t$V��豴��j j �pPj�GP��蝴���H ���^�    �O`��t��rQ�@�@�Ѓ��G`    _[��������������j�h�d�    PQ�`r3�P�D$d�    h7h�   h�rh�   �������D$�D$    ��t���,����L$d�    Y���3��L$d�    Y�������������j�h d�    PVW�`r3�P�D$d�    �|$�7��t,�t$���D$    ������N�D$�����!���V蛭�����    �L$d�    Y_^��á�rS�@U�l$��   VW��W�_dS�wx�w`UV�Ѓ��G|����   �? ��   �; ��   �wpV�_hSU���������u&�W����rhT7�@h  ��0  �Ѓ��wU���b����j j jV��  �G|��t��������G|_^][� �G|�Gx����_^][� �G|�����    ��r�6�@�@�Ѓ��    �G|_^][� �����������V������W��    �F`    �Fd    �Fh    �Fp�Fx�����F|   ^������W���d �G`t~S�\$;_xtsU�/�͉D$�����xP u����%V�������S�t$�pPj�GP�������H ���^�G|]��u�D$�_x��t�    �G`[_� �L$�Gx������t�3�[_� �̋D$��t	�Ap� �yd t�Ah� 3��y|��� ��������t$��r�t$�@�t$�@�t$�t$�t$�t$Q�Ѓ� � ��r�t$�@Q�@�Ѓ�� �������̡�rQ�@�@��Yá�r�t$�@�t$�@Q�Ѓ�� ���̡�r�@� �����̡�rV�@�t$�@�6�Ѓ��    ^��VW��跰���t$���t$�x@�t$衰���H ���_^� �����VW��臰���t$���t$�xD�t$�q����H ���_^� �����W���X����xH u3�_�V���F����ύpH�<����H �^_�����W���(����xL u3�_� V�������t$���t$�pL�t$������H ���^_� ��W�������xP u���_� V���ӯ���t$���t$�pP�t$�t$蹯���H ���^_� �������������W��蘯���xT u���_� V��胯���t$���t$�pT�q����H ���^_� �����W���X����xX u���_� V���C����t$�ύpX�5����H ���^_� ���������j�h. d�    P��$SVW�`r3�P�D$4d�    �ً|$D��tA�L$ ��������D$<    �خ���pL�D$ P���ɮ���H ��ЍL$ ��D$<���������t$H��tj��r�L$�@Q�@�С�r�L$�@V�@Q�D$H   �С�r�L$�@Q�@�D$L�����Ѓ����V����H@��t��rV�@Q�@�Ѓ��L$4d�    Y_^[��0� ��������VW�������t$�΍xH�	����H ���_^� �������������W�������x` u	� }  _� V���ѭ���t$�ύp`�í���H ���^_� �������SVW��覭���x` u� }  �$��蒭���p`�D$���P���~����H ��Ћ���r�\$�IS�I�у�;�@��rS�@�@�Ѓ�;�+���?����t$���t$�pDS�t$�(����H ���_^[� _^�����[� W�������xP u	�����_� V�������t$ ���t$ �pP�t$ �t$ �t$ �t$ �Ϭ���H ���^_� ���W��踬���xT u	�����_� V��衬���t$���t$�pT菬���H ���^_� ���W���x����xX tV���j����t$�ύpX�\����H ���^_� ���$P�t$ �D$    �D$    �D$    �D$    �D$    �D$    �  ����t,�$��t%�t$��r�t$�@�t$�@X�t$Q�Ѓ����3������������[��������������U������  V��MW�t$D��u'�E�~f� �~Ff�@�~Ff�@_^��]� �}���^�G0�V�o �Y�f(��Y�f(��Y��X'�FP�Xw�X��GH�Y��X��d$�d$ �g8(��Y��X��GP�Y��X��t$�t$(�w((��Y��D$8���G@�XO�Y��X��GX�Y��X��L$8�L$0����  �$����f �V�^((��YG0(��Y��Y�E�X�(��YGH�Y�j �X��G8�Y�j ����$   �X��GP�Y��X��G@�Y���$(  �X��GX�Y��X��D$ ��$8  �D$0��$@  �D$P��$H  �@�D$� �$��$   P��$<  P��$  P��$<  �
c  �  �f �V�^((��YG0(��YύD$8P�E�X�(��YGH���X�(��Y��Y���$�   (��YO8�Yg@�X�(��YGP�Y_X�X��X��D$��$�  �D$,��$�  �D$L��$�  �@�D$� �$��$�   P�X㍄$�  P��$D  P��$�   ��$�   �b  �|$8 �~ f�D$ �~@f�D$(�~@f�D$0��
  �O�Y�f�G0�^�X�Y��w8�(�M�X��GH�YÍ�$�   P��$  �X�(��Y��gX��$�   �O �YP�XO�X��GP�Y��_@�X�(��YF��$�   (��Y�XO�X�(��YF�X���XF��$�   �N�XN �D$�Y|$�L$ �N�XN(�X�Yt$ �Y\$ �L$�O�Y��G0�YD$ �X�Yd$�X��X��GH�YD$�X��X��GP�YD$��$�  ��$p  �O �YL$�XO�X��X���$x  �  ����$h  P��$\  �MP�j  � �\�D$`�@�\F�D$h�@�\F�D$`P��$�  P�D$x�j  �`�H�(�t$L�wW��Y�f(��Y��\�f(��\��Y��V�L$P��\��Y��\$X�^�g(�X7f(��YG0�l$`(��Yo �X��GH�Y��Xo�M�Y��X�(��YG8�Xg����$�  �X��GP�Y�P��$�  P�X��G@�Y��t$�l$��$�  �X��GX�Y���$�  �X��d$ ��$�  �  �P�H�XT$P�XL$X�D$H�X �M��$8  P��$L  P��$@  ��$H  ��$P  �%  � �\D$�D$`�@�\D$�D$h�@�\D$�D$`P��$�  P�D$x��  �~ ��O�f�^f�D$P�~@f�D$X�~@�Y�f�D$`(��YG0�X�E�M���X��GH�Y�j j ���X�(��YG8��$�   (��YO �XO�X��GP�Y��X��G@�Y���$�   �O(�Y��XO�X��GX�Y��X��@�D$� �$�D$`P��$�   P��$0  P��$�   �v]  �  �E� �D$�@�D$ P��$D  P�D$�  �@�L$��$�   ��$�   �L$P��$�   ��$�   ��$t  �  �f �V�G0�^(�Y�(��YʋEj ���X��GH�Y��X��G8�Y���$  (��Y��X��GP�Y��X��G@�Y��gX��$  (��Y��V8�X�(��Y��_0�Y��X��F0�Y��Y���$  �X?�N@�Xo�Y��G@�X��_H�Xw�Y��Y��Y��X��_8�Y��X��@�D$� �X��_P�Y��$��$  P�X��X�$�   P��$�  P��$�   ��$�   ��$�   �!\  �~�\$ �\^0�~H�L$(�~P�\$�\N8�\V@f(��Y��L$(��Y��T$�X�(��Y��X��%e  f(�W�f.ʟ��Dz
f(�f(��*��2�^��T$�L$�\$�Y��Y��Y��FH�Y��Y��Y��XV0�XN8�X^@f�T$ f�L$(f�\$0�  �F0�V8�_0�N@�Y��Y��Y��X?�Y��G@�Xw�X��_H�Xo�Y��Y��Y��X��_P�X��GX�X��Y��Y�j�X덄$T  �X�P��$X  ��$`  ��$h  �Z  �\$�D$�YFHf.�7�D$���Dz��7�L$�V0�O�f8�^@�Y�(��YG0�X�M��$�  P��$�  �X�(��YGHP�X�(��YG8��$�  (��YO �XO�X�(��YGP�X��G@�Y���$�  �O(�Y��XO�X��GX�Y��X���$�  �f  �M��\�I�\H�T$f(��Y��L$(��Y�W��X�(��Y��X���b  �d$f(�f/�vf(��f(�W�f.џ��Dz
f(�f(��'��2�^��T$�\$�Y��Y��Y�(��Y��Y��Y��^��f�T$(f�\$0f�L$8�,$�  ���\$�D$�Bb  �YD$�V0�O�f8fW 8�^@�Y��D$0f(��YG0�X�M��$�  P��$  �X�f(��YGHP�X�f(��YG8��$�  (��YO �XO�X�f(��YGP�X��G@�Y���$�  �O(�Y��XO�X��GX�Y��X���$�  �  �P�H� �XT$(�XL$0�XD$ ��$�  P��$�  ��$�  ��$�  ��$4  �MP��  �~ f�D$ �~@f�D$(�~@f�D$0��$`  WP�9
  �d$(�\$0�T$8�ȋE�I�A0�Y��YÃ��X	_^�X��AH�Y��X��A8�Y���I �Y��XI�X��AP�Y��X��A@�Y��H�I(�Y��XI�X��AX�Y��X��H��]� ��	�������)�������������� �������������U������   �}SVW�L$t�   _^[��]� �}�W�Pt�D$��tᡜr�]�@HS��   W�Ћ�r�u�Id�D$�I<�ы��D$|j/P�t����$�   jP�t����rV�@dW�@pS�Ѓ�(3���rj �@d��$�   �@��t�L$tQS��3���9t$��   �L$3�;���;���   �L$W���T$RV�uf�D$$f�D$,f�D$4f�D$<f�D$Df�D$Lf�D$Tf�D$\f�D$d�5�D$l�D$t    �Px�|$h�t��rj �@dj���   �L$ QS�Ѓ��L$F;t$�]���G��� ���_^�   [��]� ��������������U�������   �ESVW��t���_^[��]� ��r�L$�@HQ�M�@,�Ћ���   ��$�   �}W���D$����3��Pt���z  �W��L$Qf�D$f�D$f�D$$f�D$,f�D$4f�D$<f�D$Df�D$Lf�D$T�5VW���D$d�D$l    �Px�|$`��  �d$��$�   �\$��$�   �T$ �Y��Y��u�X�$�   ��r�u�L$xQ�X���$�   �Y��u�X���$�   �Y���$�   ��$�   �Y��X�$�   �X���$�   �Y��X���$�   �Y���$�   ��$�   �Y��X�$�   �X���$�   �Y��X���$�   �@d�@�Ѓ���t
�E�t$t�W��F�Rt;�������D$_^[��]� ����U������4  ��rS�@HV�@$�L$�MW�Ћ�r�M�RH�؋R<��$�   P���#�S�[f(̹   ���|$��YL$(�|$8f(��YD$@�XL$�t$P�l$h�X�f(��YD$X�X�f(��YD$H�Y���$�   f(��YL$0�Y��XL$�Xd$ �X�f(��YD$`�X��S(�Y��X��X��[ ��$�   f(��YD$@��$�   �cf(��YL$(�X�f(��YD$X�X�f(��YD$H�Y���$�   f(��YL$0�Y��X�f(��YD$`�X��Y��X��X���$�   ��$�   �[8�c0�S@f(��YL$(f(��YD$@��r�uj �X�f(��YD$\V�X�f(��YD$P�Y���$   f(��YL$8�Y��X�f(��YD$h�X��[P�Y��X�f(��YD$H�X��SX��$  ��$  �cHf(��YL$0Ǆ$�       �X�f(��YD$`�X�f(��YD$P�Y���$  f(��YL$8�Y��X�f(��YD$h�X��Y��X�W�f�D$xfք$�   fք$�   fք$�   fք$�   fք$�   fք$�   fք$�   fք$�   �5�X���$�   �@@��$   �@8��$(  �Ћ}����L$pQWV���Rx�u�\$��$�   �3P�u��$4  P��$�   �n����~ �L$pQ����W�uf��~@f�A�~@f�A���V|_^�   [��]� �3�� �����������3�� ������������ �������������3�� ����������̸   �$ ��������� �������������3�� ������������ �������������3�� ������������ ��������������$ ������������̡�r�L$�@��   �@<�Ѕ�t#j ��$8  ��$,  � �������u��   �Sh   �D$j P��V  ��$<  j ��$L  �D$��$T  S��$P  P�   ��$�   ����E���$�   ��$�   �� ��E���$�   ��$�   �À��E���$�   ��$�   ����E�h   ��$�   �D$,P��$X  Ǆ$�   ���$X  j�	g����8[��   ���������������V�t$W�t$ �|$�t$V�t$�t$$W���������   Ǉ�   �Ǉ�   �Ǉ�   �Ǉ�   ��Ǉ�   �Ǉ�   ��Ǉ�   �_^��������������U�������   VW�M�qX�I8�y(�A@�YAP�Y�f(��YQP�D$X�L$H�\��A �D$`�Y�f(��T$8�Q �YQ@�\��D$h(��YA8�T$ �L$0�D$(��Q0�\��A�Y��Y�W��|$(�\$@�X��AH�Y��d$P�X���2f.џ��DzD�Ef�f�@f�H0f�HHf�Hf�H f�@8f�HPf�Hf�H(f�H@f�@X_^��]��^��y�D$�A(��Y�(��Yq@(��Ya8�(��YYP(��Yy �\��d$(��\��d$h�YA0�\d$8�YIH�\t$�\��i�X��D$X�\D$H�Y��Y��Y��Y��X��YL$�L$p�I�YL$((��\��\��YAH�Yy0�X��X��\$�Y��D$x�D$�\D$ �Y��QH(��YI@�X��D$0�Y��X��y0��$�   �D$@�Y��Y���$�   �D$P�Y���$�   ��$�   (��YAX�\�(��YA(�Y���$�   (��YIX�\��Y���$�   (��YI((��YA@�E�t$p���\�(��YA8�YT$`�Y���$�   (��YIP�Y|$`�\�(��Yi8�YAP�Y��\��\й   ��$�   �Y��Y���$�   ��$�   �_^��]����U����QV�u�V��^(��Y��Y��X�(��Y��X��JS  f(�W�f.џ��D�Ez��H�H^��]���2�^���Y���N�Y��H�N�Y�^�H��]Ë�`D��`H��`L��`P��`T��`X��`\��``��`d��`h��`l��`p�������������L$f/�2r��7���7f/�r��7�(��bR  �D$�D$�̡�r���@h�t$ �@0Q�L$Q�ЋL$(�~ f��~@f�A�~@f�A����$� �������������̡�r���@h�t$ �@8Q�L$Q�ЋL$(�~ f��~@f�A�~@f�A����$� �������������̡�r���@h�t$ �@,Q�L$Q�ЋL$(�~ f��~@f�A�~@f�A����$� ��������������h�rjh�f �<  ����t	�@��t�����������������j�hX d�    PQV�`r3�P�D$d�    h�rjh�f �D$     �5<  ������t9�~ t3�t$L�D$$�t$L�t$L�t$L�t$L����P�Ð���t$L�F�Ѓ�4�������L$ �D$���������ƋL$d�    Y^���������������h�rjh�f �;  ����t	�@��t��3��������������h�rjh�f �;  ����t�x t�@��3������������h�r�t$h�f �M;  �����������̋D$HV����   �$����   ^á�r@��r��uX�t$������=�2  }�����^Ët$��t�h8jmh�rj�n�������t	��� ����3���r��tV�������   ^��t$�t$�'n���������H^�^��m����ru.��m��袶���5�r��t��豏��V�+�������r    �   ^Ã��^Ë�ݫf�l�֫��L����������L$u�D$��r�D$��r�   � �� �h6V���.�vf(�fT 9f/�f(�fT 9�T$�L$�L$�-  f/��#  ��8f/�vFf/�v@�,��,���   ��$    ������ʅ�u�fn�����^��^��.�v^�� �f/�v(��(���8�^��%�2f/�v4(��Y��Y��Y��D$(��Y��.�v(��L$�L$f/�v(��D$�D$�f��D$�D$�M  �\$�D$f/�8�L$�L$�D$�D$s���^���F�^��F^�� �W����2�F^�� �����������������D$��8f/�V��w��8f/�v(��Y(5���X�8�D$�D$�$��K  �(5������F�������^� ���̃��L$�T$3�W�f/�fT 9�X�8��3�f/�V����3��L$�D$;������$�L$�gK  ��D$ fT 9�D$ �X�8�D$ �D$ �$�7K  ��2�\$ �D$ ��f/��Fv'��rhX8�@j��0  ����2���F�|$ u�fW 8���������^��� ������������D$��2f/�V���Fv'��rh�8�@j,��0  ����2���F^� ���������U�����M��2��<f/�V��v'��rh�8�@j5��0  ����2���M��Y����D$8�D$8�$�J  �\$8�F�$��I  �D$8�\$@�^D$@�D$@�D$@�$��I  ��E�$��I  ���^�������^��]� ����������̡�rQ���   �@X�Ћȃ���u� ��r�t$�@|�t$�@Q�Ѓ�� ������̡�rQ���   �@X�Ћȃ���u� ��r�t$�@|�t$�@8Q�Ѓ�� ������̋T$V��j ���rj �@j �@R�Ѓ��F��^� ������̡�rV�@j �@j ��j �6�Ѓ��F^�V��N��u3�^� ��rQ�t$�@�t$�@�6�Ѓ��F�   ^� ��������̋L$��`������̋L$��`�������V��hP��9�F    ��rV�@Ph0�� h ��Ѓ��F��^����������̃y �9u��r�q�@P�@��Y��̋I��u3�� ��rj �t$�@P�t$�@Q�Ѓ�� �����̋I��t��r�t$�@PQ�@�Ѓ�� ̋I��t��r�t$�@PQ�@�Ѓ�� ��    �A    ���V����t&��rQ�@P�@L�С�r�6�@P�@<�Ѓ��    ^����������������SUVW�����t��rQ�@P�@<�Ѓ��    �G    �\$�l$hP�S�o��rh0��@Ph ��@8U�t$(�Ѓ�3����~D���x u�@   ��r�HP���p�A�Ѓ���rV�@P�7�@@�Ћ�F���A;�|�3�9_^]��[� �������������t$�D$�t$�p�,���� ���������SVW��3�9w~>�\$��rV�@P�7�@@�ЋЃ���t,��rj �APS�@jR�Ѓ���tF;w|�_^�   [� ��r�7�@P�@L�Ѓ�3�_^[� ̡�r�1�@P�@D�Ѓ��������������̡�r�1�@P�@H��Y���������������̡�r�1�@P�@L��Y���������������̡�r�@P�@P����̡�r�@P�@T����̡�r�@P���   �࡜r�@P���   ���L$��`�������V��~ �9u��r�v�@P�@�Ѓ��D$t	V�1}������^� ��������3��������������̡�rQ�@D�@$�Ѓ���������������̡�rj �@D�t$� �Ѓ�����������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@D�@�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�r�@D� �����̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�r�t$�@Dh2  � �Ѓ��������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�rj �@D�t$� �Ѓ�����������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�r�t$�@Dh'  � �Ѓ��������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�r�t$�@DhO  � �Ѓ��������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�r���@XQ� �L$Q�ЋL$$�~ f��~@f�A�~@f�A���� � ��̡�r���@XQ�@�L$Q�ЋL$$�~ f��~@f�A�~@f�A���� � �̡�r���@XQ�@�L$Q�ЋL$$�~ f��~@f�A�~@f�A���� � �̡�r��`�@XV�@WQ�L$Q�Ћ��D$t���   ���_^��`� �������������̡�r�t$�@XQ�@�Ѓ�� �������̡�r�t$�@XQ�@�Ѓ�� �������̡�r�t$�@XQ�@�Ѓ�� �������̡�r�t$�@XQ�@�Ѓ�� �������̡�r�t$�@XQ�@$�Ѓ�� �������̡�r�t$�@XQ�@ �Ѓ�� �������̡�rj �@Dh�  � �Ѓ����������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@D�@(�Ѓ���������������̡�rQ�@D�@�Ѓ���������������̡�r�t$�@D�t$�@Q�Ѓ�� ���̡�rj �@Dh:  � �Ѓ����������̡�rV�@@�t$�@�6�Ѓ��    ^�̃���r�$    �D$    ���   �$�@Rj�����#D$��������������̡�rj �@Dh�F � �Ѓ����������̡�rV�@@�t$�@�6�Ѓ��    ^�̋D$����u��� �D$��r�$    ���   �$�@Rj������؃�� �̡�rj �@Dh�_ � �Ѓ����������̡�rV�@@�t$�@�6�Ѓ��    ^�̡�rQ�@\�@�Ѓ���������������̡�rQ�@\�@�Ѓ���������������̡�r�t$�@\Q�@�Ѓ�� �������̡�r�t$�@\�t$�@Q�Ѓ�� ���̡�r�t$�@\Q�@�Ѓ�� �������̡�rQ�@\�@�Ѓ���������������̡�r�t$�@\Q�@ �Ѓ�� �������̡�r�t$�@\�t$�@$Q�Ѓ�� �����t$��r�t$�@\�t$�@(Q�Ѓ�� ��r�t$�@\Q�@0�Ѓ�� �������̡�r�t$�@\Q�@@�Ѓ�� �������̡�r�t$�@\Q�@D�Ѓ�� �������̡�r�t$�@\Q�@H�Ѓ�� �������̡�rQ�@\�@4�Ѓ���������������̡�r�t$�@\�t$�@8Q�Ѓ�� ���̡�r�t$�@\Q�@<�Ѓ�� ��������QSUVW�|$��j ���<�����rU�@\�@�Ѓ���S���!���3���~B�	��$    ����r�L$�@\Q�@(�L$QVU�Ѓ����t$�����t$���ޒ��F;�|�_^][Y� ̃�S�\$W�D$��P�������|$ ��   ��rW�@\�@�Ѓ��D$P��������D$��taV3���~L���D$P��褔���D$P��蘔���L$;L$!��rQ�@\W�@�ЋL$$A���L$;L$~�F;t$|�^_�   [��� _�   [��� ����������̡�r�@\� �����̡�rV�@\�t$�@�6�Ѓ��    ^�̃�S�\$$�щT$���.  �L$(U��V��EW�}��C���|$,��D$,���މt$$���l$ �|$�D$�t$��l$ �|$�t$���~t$$M+��l$ �t$�|$�A�P����t+��D�J�R��Nu�L$4�D$K�\$0����   �T$�t$+��D$�<m    ;����w���t$,;�}��SV�����yG��\$0�L$V�U��L$4�T$���D$�I����F��م�t+�L(�P�@��(Ku�L$4�\$0�T$�;�~��D$����_^][��� ���̃�S�\$(�L$�L$,U�����l$���D  V�t$,W����G�|$�G�����C���D$0���ۉ\$(�\$4�t$�D$�t$ ��I �l$$�|$�t$�d$ ��~�T$(T$ O+�|$�t$�L�P�����t/�|$+���$    �Jf�D�Rf�f�Nu�L$8�|$�D$K�\$4����   +��D$�T$�t$ �;����w���t$0;�}��SV�����yG��\$4�L$V�U��L$8���D$�<����L$$�F��م�t+��Pf�L(�@f�f�(Ku�\$4�L$8�T$�;�~��D$�����_^][��� �̃�S�\$(�L$�L$,U�����l$���<  V�t$,W����G�|$�G�����C���D$0���ۉ\$(�\$4�t$�D$�t$ ����l$$�|$�t$�d$ ��~�T$(T$ O+�|$�t$�H�P�����t+�|$+���$    �D�J�R��Nu�L$8�|$�D$K�\$4����   +��D$�T$�t$ �;����w���t$0;�}��SV�����yG��\$4�L$V�U��L$8���D$�@����L$$�F��م�t+L(�P�@��(Ku�\$4�L$8�T$�;�~��D$����_^][��� ��������̋T$�T$������3������� ������������������Q�D$SW�L$��t+�\$��t#�|$��t�|$ t�SP���u_��[Y� y_3�[Y� U�   OV;�|1���L$�4/������\$$\$S�t$���ty�~���n;�~�^]_3�[Y� ��~-�l$$���|$$��|$���L$��W�t$N���u�߅��^]_��[Y� �����������̋D$SUW�����   �\$����   �|$����   �|$ ��   �U SP���u_]��[� y�D$ _]�     3�[� �   VO3��L$;�|:�d$ �E �4�����\$ \$��S�t$���t*y	�L$�~���N�L$;�~ʅ��D$$~F�0^_]3�[� ��~2�D$ ���|$ ��|$�D$$��E W�t$��N���u
�D$$�߅��^_]��[� �D$ _]� ����3�[� ������    �A    �A    �A    �����V��V��m���FP��m�����F    �F    ^������������S�\$V��W�~�    �    �F    �F    �CV;C��   �m��W�m���F    �F    ��rh$9�@jI���   j�Ѓ������   ��rhP9�@jN���   j�Ѓ����uV�6m������_^[� ��F   �F   ����C�A��C�A�_�    ��^[� ��l��W��l���F    �F    ��rh$9�@jI���   j�Ѓ����tZ��rhP9�@jN���   j�Ѓ�����Z�����F   �F   ����C�A��C�A��C�A��    _��^[� ����������V�t$���    �F    �F    �F    �  ��^� ���V�t$���  ��^� ��������������SUV��V��k���nU��k���\$���F    �F    ��t(��rh$9�H��    jIP���   �Ѓ����u^]3�[� W�|$��t;��rhP9�H��    jNP���   �Ѓ��E ��uV�kk����3�_^][� �~_�^^]�   [� �������������V��V�7k���FP�.k�����F    �F    ^������������SV��WV�k���^S��j���|$���F    �F    ����   �? ��   �W����   ��rh|9�H��    jlP���  �Ѓ����t<� t>�W��t7��rh�9�H��    jqP���  �Ѓ����u���'���_^3�[� �G��F�G�FQ��PQ�7�4�������t�FQ��PQ�w�����_^�   [� ������������SUV��WV�j���~W��i�����|$ �F    �F    �  �\$����   ��rh�9�@��    ���  h�   Q�Ѓ����tB�l$ ��tL�T$��tD��rh :�H��    h�   P���  �Ѓ����u���&���_^]3�[� �D$�F�,�F   ��rh,:�@h�   ���  j�Ѓ����t���^��t��    ��tQ�t$ P��.  ����t ��FQ��PQU��}�����   _^][� ��_^]�   [� ���    �A    �A    �A    �����U������   �U��V�HWW�3��<��D$�|$@�L$}
��_^��]� ����  �0�U�f(ύ@�F�~ʍ@f(��D��,��t��\D��D$�\t��8�L$(�|$ �T$�\$0�\��D$8����   ��������f(ƍ@f(��$��T��\T��\��\��\\����Y��Y��Y��Y��\�f(��Y��Y��XL$(�\�f��\$0�\��L$(�Xl$�Xt$ �l$f�f(��D$ f�O�f����T$W��(��YL$(�YD$ �}f�?�X�f(��Y�f�f��X���-  �T$(�\$ f(�W�f.͟��Dz�L$f(�f(�f(��&��2�^��L$f(�f(��Y��Y��Y�f�gH�% 9fT�fT�f/�f�wPf�GX��   f(�fT�f/���   �GH�WX�gP(��Y�(��Y��\��Y��\�f�_�\�f�O f�g(�OX�P�Y(�W�gH(��YG (��YWP�\�(��YG(�Yg �Y�f�0�\��\�f�_8f�g@�)  �WPfT�f/��_X��   �OH�Y�f(��Y��\��\��Y�f�Gf�_ �\�f�O(�(�G �YGX�YP�O�wH(��Y_X�YOP�\�f(��YG(�Yw f�0�\��\�f�_8f�w@�   f(��Y�(��Y��\��GH�Y�f�O0�\��\�f�_8f�G@�oP�X�Y8�OH�w0(��YG@(��Y_@�YO8�\�(��YGX�Y�f��\��\�f�_ f�w(�D$`WP������U���D$�   ���W�3�3Ʌ�~w��r]�p��W�W�%  �yH���@��+���    �o���f���oD��f��;�|�f��fo�fs�f��fo�fs�f��f~ϋt$;�}�F<�A;�|���t$�M��u�A0�D$(���q �@�D$    ���d��\��Y�f(��YI�D$(�Y��X	�D��Xq�@�X��AH�Y��X��A8�Y��L$ �I(�X��AP�Y��Y��T��X��A@�XI�Y��$��X��AX�Y�(��YY�X�(��YA0�Xf�L$X�L��D$�X�(��YAH�@���X�(��YA8�YQ@�\$(��YY �Ya(�D$�XY�Xa�X�(��YAP�YIX�X��X��X��\$0f�d$8���  3�������|$�D$(׋��@�,��T��L�f(��Ya(��YA0�X!f(��YY �Yi(�X��XY(��YAH�Xi�D$@�X�(��YA8�YQ@�D$�X�(��YAP�YIX�X��T$0�X�(��X�f(��\��\��\�f�\$0�YL$�YD$ �Y��X��~D$�D$ �~D$8f�D$X�X�f�f�d$f�l$8�X�;D$������|$@�D$@_^��]� �����������̋�����������T$�   @t������@��wm�$����D$� ����D$� ���� �
�D$��D$�J�� �J�D$��D$�J�� �J�D$��D$�J�� �J�D$��D$�
�� �I ����������S��V�����%���W��   @t�����ʃ��|$;�t�����t�t$�����t��t$;�t>�����t6�΁����Eǃ��t����   �_�^�[� ��   ���Ё�   @�_^[� ���U�������AW�SVf(�f(�f(�W�L$�\$�T$ �D$���L  �9�u������Ш�)  ���������U��Z�@�[�<��l��\<��\l�;Zuc�\��B�\\��@�d��\d��T��\T��4��\4�f(��Y�f(��Y��Y��\�f(��Y��\��Xd$(��d�d��B�\d��@�B�@�T��\��\\��\T��4��\4�f(�f(��Y��Y��Y��\�f(��Y��\��X\$�XL$�Y��Y��\$�L$�\��Xt$ (��T$ ���L$�����f(��Y�f(��Y��X�f(��Y��X��%  f(�W�f.П��D�Ez� �@�@_^[��]� ��2�^�_^[(��YD$� (��YD$�@�D$�Y��@��]� ���������U������<�05�585�AS3�Vf�f�f�f�W�D$�L$�|$ �t$(�l$0�d$8�T$@�D$���4  ��u��    ������Ш��  ���������M��@��ts��f/�v
f(��D$�\�f/�v
f(��L$�\�f/�v
f(��|$ f/�v
f(��t$(�T�f/�v
f(��l$0f/�vPf(��D�~4��~l��~d�f�f�f�   �t$(�l$0�D$�L$�|$ �T$@�d$8�A�@��ts��f/�v
f(��D$�\�f/�v
f(��L$�\�f/�v
f(��|$ f/�v
f(��t$(�T�f/�v
f(��l$0f/�vPf(��D�~4��~l��~d�f�f�f�   �t$(�l$0�D$�L$�|$ �T$@�d$8�y���ts��f/�v
f(��D$�\�f/�v
f(��L$�\�f/�v
f(��|$ f/�v
f(��t$(�T�f/�v
f(��l$0f/�vPf(��D�~4��~l��~d�f�f�f�   �t$(�l$0�D$�L$�|$ �T$@�d$8�A;�t8�@�L$��P�E  �T$@�d$8�l$0�t$(�|$ �L$�D$���L$�@�����te�Ef(��X�f(��X���8f(��X��Y��Y��Y�f�f�Pf�H�\0�\h�\`�Ef�0f�hf�`_^[��]� �EW�f� f�@f�@�E_f� ^f�@f�@[��]� ��������̋Q3���|�	��t��~�    t@��Ju��3����������̋QV�t$��;�}�	���    u@��;�|����^� +�@^� ���������������VW�|$���x*���t$�v3Ʌ�~��I ���%���;�tA��;�|�_���^� _��^� �����������SV�q2ۅ�~;�W�|$�
����%���;�u��   @u�����t	�   ���3�
؃�Nu�_��^��[� V�q3҅�~�	�d$ ��   @u	�����tB��Nu��^�����V�q3҅�~�	�d$ ����ШtB��Nu��^�����������QV��3�9N~��I �A�d�����;N|��N��~gSU3�W�   �T$����x;���������;�},�I ����<����������;�u��   ��@;F|ۋT$�NE���E��T$;�|�_][^Y����������������h�rjh_� �O
  ����uË@����V�t$�> t1h�rjh_� �%
  ����t��L$�@�L$Q�Ѓ��    ^����Vh�rjh_� ����	  ����t�@��t�t$����^� 3�^� ������������Vh�rjh_� ���	  ����t�@��t�t$����^� 3�^� ������������Vh�rjh_� ���l	  ����t�@��t�t$���t$�t$��^� 3�^� ����Vh�rjh_� ���,	  ����t�@��t�t$����^� 3�^� ������������Vh�rj h_� ����  ����t�@ ��t�t$����^� 3�^� ������������Vh�rj$h_� ���  ����t�@$��t�t$����^� 2�^� ������������Vh�rj(h_� ���l  ����t�@(��t��^��3�^������Vh�rj,h_� ���<  ����t�@,��t��^��3�^������Vh�rj0h_� ���  ����t�@0��t�t$����^� 3�^� ������������Vh�rj4h_� ����  ����t�@4��t�t$���t$��^� ���^� �������Vh�rj8h_� ���  ����t�@8��t��^��3�^������Vh�rj<h_� ���\  ����t�@<��t�t$����^� ��Vh�rj@h_� ���,  ����t�@@��t�t$����^� ��Vh�rjDh_� ����  ����t�@D��t�t$����^� 3�^� ������������Vh�rjHh_� ���  ����t�@H��t�t$����^� ��Vh�rjLh_� ���  ����t�@L��t��^��3�^������Vh�rjPh_� ���\  ����t�@P��t��^��3�^������Vh�rjTh_� ���,  ����t�@T��t��^��^��������Vh�rjXh_� ����  ����t�@X��t��^��^��������Vh�rj\h_� ����  ����t�@\��t��^��^��������Vh�rj`h_� ���  ����t�@`��t�t$���t$��^� 3�^� ��������Vh�rjdh_� ���\  ����t�@d��t�t$���t$��^� 3�^� ��������Vh�rjhh_� ���  ����t�@h��t�t$���t$�t$�t$�t$��^� ��Vh�rjlh_� ����  ����t�@l��t�t$���t$�t$��^� 3�^� ����Vh�rjph_� ���  ����t�@p��t�t$���t$��^� 3�^� ��������Vh�rjth_� ���\  ����t�@t��t�t$���t$��^� 3�^� ��������Vh�rjxh_� ���  ����t�@x��t�t$���t$��^� 3�^� ��������Vh�rj|h_� ����  ����t�@|��t�t$����^� 3�^� ������������Vh�rh�   h_� ���  ����t���   ��t�t$���t$��^� 3�^� ��Vh�rh�   h_� ���Y  ����t*���   ��t �t$���t$�t$�t$�t$�t$��^� ���^� �Vh�rh�   h_� ���	  ����t*���   ��t �t$���t$�t$�t$�t$�t$��^� ���^� �Vh�rh�   h_� ���  ����t"���   ��t�t$���t$�t$�t$��^� 3�^� ����������Vh�rh�   h_� ���i  ����t���   ��t�t$����^� 3�^� ������Vh�rh�   h_� ���)  ����t���   ��t�t$����^� ������������Vh�rh�   h_� ����  ����t���   ��t�t$���t$��^� 3�^� ��Vh�rh�   h_� ���  ����t���   ��t�t$���t$�t$��^� 3�^� �������������̃��L$�T$�D$�R�X�A�\B�\��\Y�Y �Y�Y�X��X��$�$�������h�r�t$h_� �  �����������̃y0 �D$tq��f/�v�	�H�Af/�v�I�H�Af/�v�I� f/Av�A�@f/A v�A �@f/A(vI�A(� �~ f�A�~@f�A �~@f�A(�~Af��~A f�A�~A(f�A�A0   � ̋L$�D$Q��D$j�t$�A�S-�������������������̸   �����������V�t$��t���u7j�t$�6-������u3�^Ë���,���ȅ�t��t��D$3�;AOʋ�^��������̋ыB��:��t!�J��t�H�J�B�A�B    �B    ���������������̋T$�B�A�J�A�Q�H� ������̋T$�B�A�J�A�Q�H� ������̋ыB��t!�J��t�H�J�B�A�B    �B    ��������:�A�:�A    �A    �Q�A� �:�@    �@    �A�A    �A    �Q�A    ����������������j�h� d�    PQV�`r3�P�D$d�    ��t$��:�D$   �  �N�F�:��t!�F��t�A�N�F�A�F    �F    �N�F�:��t!�F��t�A�N�F�A�F    �F    �L$d�    Y^��������̋A��3�V;�t ��t�t$��B;�t�@��t
�x t��u�3�^� ������������̋A�T$�B�A�B�A�P�Q� ���̋T$�A�B�A�B�A�P�Q� ���̍A�A�A�A    �A�A    ������SW���O�_;�t!��tV�q��t�~ u3��j��΅�u�^�G�_�G    �G�G    _[�������̋A��;�tE��tAV��H��t
�y t���3��P��t��t�J�P�H�J�@    �@    �ƅ�u�^ËQV�A3�;�t��t�RF��t
�z t��u��^����������VW���wV��:�}J�����G    �G    _�    ^����S�\$V��F;�~��x�N�D$��^�   [� ^3�[� }hW�~9~uI��u�~��F��t�����t?��rhX:�Hj8��    P�v��  �Ѓ���t�F�~�N�F��    �F9^|�_�F;Fu����  ���x����V�N�D$���F^�   [� ������̋T$V���x)�F;�}"�L$��x;�};�t�F�4��������^� �������̋T$V�t$W��;�}N��x.�G;�}'��x#;�};�t�GS��R�k  ��t	VS����   [_^� �������̃��D$j�q�D$�:�q�L$�D$������� �����̃��D$j�q�D$�:�q�L$�t$�D$������� ��VW���O�q���x6;�}2�G����t*��x&;�}"�w;�}��I �O��F�J�
;w|�_^�3�_^��������V��F;Fu�p  ��u^� �V�N�D$���F�   ^� ���������������V��W�F�|$;�O�3Ʌ�H�;Fu���  ��u_^� �F;�~�N��H�J��
;���N�D$���F_�   ^� �����̋T$V���x/�F;�}(H�F;�}��    �F��B�A�;V|�   ^� 3�^� V��3ҋNW��~�F�|$98tB��;�|�����x);�}%�A��F;�}�F��B�A�;V|�_�   ^� _3�^� ��������̋Q3�V��~�I�t$91t@��;�|���^� �������������A    ���������VW���wV��F�����G    �G    _�    ^����������QSUV�t$W���nU�|$�F���E     �F    �F    �G�F�G3ۃ��F9_~u�G�~���D$9~uI��u�~��F��t�����tV��rhX:�Hj8��    P�u ��  �Ѓ���t-�E �~�N�E �T$�|$���FC;_|�_^]�   [Y� _^]3�[Y� �V��W�~��u�~��F��t�����u_3�^á�rhX:�Hj8��    P�v��  �Ѓ���t҉~�F_�   ^����VW���wV��:�]E�����D$�    �G    �G    t	W��B������_^� ���������������V���h����D$t	V�B������^� ��V��F��:��t!�N��t�H�N�F�A�F    �F    �D$t	V�rB������^� ����������t$�A�t$�Ѓ�� ������������̡�r�@d�@P����̋L$�9 t��r�L$�@d�@T���������t$��r�t$�@h�t$� �t$Q�Ѓ�� ��������������t$��r�t$�@h�t$���   �t$Q�Ѓ�� ����������t$��r�t$�@h�t$�@Q�Ѓ�� �t$��r�t$�@h�t$�@ �t$�t$Q�Ѓ�� ���������t$��r�D$�@h�����   �$Q�Ѓ�� ��������t$��r�D$�@h�����   �$Q�Ѓ�� ������̡�r�t$�@h�t$���   Q�Ѓ�� ̡�r�t$�@h�t$���   Q�Ѓ�� ��D$��r���@h�t$<���   �t$<���D$�D$@�$�t$<�t$<Q�L$$Q�ЋL$D�~ f��~@f�A�~@f�A����@�$ ������D$��r���@h�t$8���   ���D$�D$<�$�t$8�t$8Q�L$ Q�ЋL$@�~ f��~@f�A�~@f�A����<�  ���������j�h� d�    P��VW�`r3�P�D$$d�    ���D$    �|$4�    �G    �D$8�D$�D$P�L$�D$0    �D$   �D$     �D$$    ��q��j W�D$P���D$8   ��m���L$�D$, �Us���ǋL$$d�    Y_^��$� ����������������t$��r�t$�@h�t$���   �t$Q�Ѓ�� ��������̡�r�t$�@hQ���   �Ѓ�� ����̡�r�@h�@X����̋L$�9 t��r�L$�@h�@\�������̡�r�@h���   ���t$��r�t$�@h�t$�@`�t$�t$�t$�t$Q�Ѓ� � �t$��r�t$�@h�t$�@d�t$�t$�t$�t$Q�Ѓ� � ��r�t$�@h�t$�@hQ�Ѓ�� ���̡�r�t$�@h�t$�@lQ�Ѓ�� ���̡�r�t$�@h�t$�@pQ�Ѓ�� �����t$��r�t$�@h�t$���   �t$�t$�t$�t$Q�Ѓ� � ��������������t$��r�t$�@h�t$���   �t$�t$�t$�t$Q�Ѓ� � ��������������t$��r�t$�@h�t$���   �t$�t$�t$�t$Q�Ѓ� � ��������������t$��r�t$�@h�t$���   �t$�t$Q�Ѓ�� ������t$��r�t$�@h�t$���   �t$Q�Ѓ�� ����������t$��r�t$�@h�t$�@tQ�Ѓ�� ��r�t$�@hQ�@x�Ѓ�� �������̡�r�@h���   ���t$��r�t$�@h�t$�@|Q�Ѓ�� �t$�D$��r���@h�D$�D$(���   �D$�D$ �$Q�Ѓ� � ;`ru���K  �%�0U���EV��t%Wh���~��7jV�  �EtW�;��Y��_���  �EtV�;��Y��^]� Vh�   �80Y��V�0��u��u��u3�@^Ã& �  h���V  �$* �J  Y3�^�U��QQ�} SVW�)  ��r���  H��rd�   3��P�}���u�;�t3�������u���E�   �=�utj�  Y�  �5�u�0���u����   �5�u�0�؉u�]��;�r\9;t�W�09t��3�0W���0����5�u�50���5�u�E��֋M�9Mu�u9Et���M�u�E��띃��tV��0YW�0��u��u��u�=�u9}���   3���   3��   �}��   d�   3��P����u�;�t3�������u��3�F9=�uj_t	j�  �5h�0h�0��u   �  YY��u�h�0h�0�  Y�=�uY��u3���=�u th�u�  Y��t�uW�u��u��r3�@_^[�� U��}u��  �u�u�u�   ��]� jh�b�  3�@���u�3ۉ]��}�=pr�E���u9=�r��   ;�t��u8��:��t�uW�u�Ћ��u����   �uW�u�������u����   �uW�u�ʲ�����u��u.��u*�uS�u谲���uS�u�@�����:��t	�uS�u�Ѕ�t��uK�uW�u�������#��u�t4��:��t+�uW�u�Ћ���M�� �E�QP�c  YYËe�3ۋ�u�]��E������   ����  Ëu��pr�������%�0�%�0�%|0�%x0�=�u t3��Vjj �P0YY��V�0��u��u��ujX^Ã& 3�^�jh�b�(  �5�u�50�։E���u�u�X0Y�ej�{  Y�e� �5�u�։E��5�u�։E��E�P�E�P�u�50��P�S  �����}��u��֣�u�u��֣�u�E������   ����  Ë}�j�  Y�U���u�P��������YH]��%t0�%L0�%$0�%(0U���0j��u��  �u��  �=�u YYuj��  Yh	 ���  Y]�U���$  j��  ��tjY�)��s��s��s��s�5�s�=�sf��sf��sf��sf��sf�%�sf�-�s���s�E ��s�E��s�E��s�������s  ��s��r��r	 ���r   ��r   jXk� ǀ�r   jXk� �`r�L�jX�� �dr�L�h�:�������jh�b�   �e� �]�Ë}�ǋu��u�e� O�}x+�u���U��3�@�E��E������   �!  � �}�]�u�E��u�uWSV�   �jhc�  �e� �Mx:�M+M�M�U��E�E�E� �E��E��8csm�t�E�    �E���  �e��E������  � ��%,0�%00�%40������������U��ES�H<�V�A�Y��3��W��t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�h8ch� d�    P��SVW�`r1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��E�MZ  f9t3�]ËH<�3��9PE  u�  f9Q��]�U����`r�e� �e� VW�N�@��  ��;�t��t	�Уdr�f�E�P�0�E�3E�E�� 01E��01E��E�P�0�M�3M�E�3M�3�;�u�O�@����u��G  ��ȉ`r�щdr_^��VW�<C�<C����t�Ѓ�;�r�_^���VW�DC�DC����t�Ѓ�;�r�_^���%<0�%@0h�u�   Y�����������h� d�5    �D$�l$�l$+�SVW�`r1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�U���u�u�u�uh��h`r�5   ��]��%H0�%�0�%T0�%\0�%`0�%d0�%h0�%l0�%p0�%0�������̍M��^���M��0;���M������T$�B��J�3�������C�����������������h�0jnh�r�E�P�+5����ÍM�����M��i���T$�B��J�3��G����`C�L���������������h�0h�   h�r�E�P��4����ÍM��L���M��Ti���T$�B��J�3��������C�������������̋E���   �e���M���ËT$�B܋J�3������@D�����M������M������M���h���T$�B؋J�3������D������������̋M������T$�B��J�3��X����F�]����������������h�2h�   h�r�E�P��3����ËM�����T$�B��J�3������tD����̍M�8���M�� d���M���c���T$�B�J�3��������E�����������������̍M������T$�B̋J�3�������E����������������̍M�����M������M���8���M���8���M�����T$�B��J�3��X�����D�]���������������̍M��[���M��p���M��h���M�����M��(c���M�� c���M��H���M��@���M��8���M��p���M���b���M���b���T$�B��J�3�������E���������̍M������M������T$�B؋J�3�������D��������̍M��8���Eԃ�t�e���M��7��ËT$�B��J�3��c����@F�h����������̋M�����T$�B��J�3��8�����J�=����M��e���T$�B��J�3�������J�����M��B���T$�B��J�3��������J������M�����T$�B��J�3�������tJ������M������T$�B��J�3������PJ�����M������E����   �e���M����ËT$�B�J�3��p����,J�u����M���6���M����Eԃ��   �e���M�6��ÍM��t���T$�B؋J�3��$����J�)����M��6���M�I���Eԃ��   �e���M�q6��ÍM��(���T$�B؋J�3��������I������M��E6���Eԃ��   �e���M����ÍM������T$�B��J�3�������I�����M�����E����   �e���M��5��ËT$�B��J�3��X�����I�]����M�����T$�B�J�3��5����xI�:����M��b���T$�B�J�3������TI�����M��?���T$�B�J�3�������0I������M��\5���M����Eԃ��   �e���M�<5��ÍM������T$�B؋J�3������I�����M��5���M�����Eԃ��   �e���M��4��ÍM�����T$�B؋J�3��W�����H�\����M�����E����   �e���M�l��ËT$�B�J�3�������H� ����M��4���M��@���T$�B��J�3��������H������M��]4���M����Eԃ��   �e���M�=4��ÍM���
���T$�B؋J�3������|H�����M��4���M��
���Eԃ��   �e���M��3��ÍM��
���T$�B؋J�3��X����XH�]����E����   �e���M��3��ÍM��l
���E����   �e���M��3��ËM�K
���E����   �e���M�s3��ÍM��*
���M��"
���T$�B��J�3�������4H������M��?3���M��	���Eԃ��   �e���M�3��ÍM���	���T$�B؋J�3������H�����M��	���E����   �e���M�	��ËT$�B�J�3��J�����G�O�����������������̍�h����2����X����Z	���M��2���M��2���M��2���M��z2���T$��\�����X���3�������<K�������������̍M��(U���T$�BЋJ�3�������Q�����M��U���T$�B�J�3�������Q�����E����   �e���M�����ÍM������T$�B�J�3��Y�����Q�^����M��T���M������T$�BԋJ�3��.�����Q�3����M��{T���M��c����T$�B��J�3������\Q�����M��PT���M��8����T$�B��J�3�������8Q������M��%T���M������T$�B؋J�3������Q�����M������T$�B�J�3�������P�����M�����T$�B�J�3��g�����P�l����M�����M�����T$�B܋J�3��<�����P�A����M��0���M��0���M��Y���T$�B��J�3��	�����P�����M��6���T$�B�J�3�������`P������M��S0���T$�B��J�3�������<P������M��S���M�������M�������M�������T$�B؋J�3������P�����M���R���T$�B�J�3��e�����O�j����M��R���T$�B�J�3��B�����O�G����M��R���T$�B�J�3�������O�$����M��lR���M��T����T$�B؋J�3��������O������M��AR���M��)����T$�B؋J�3�������dO������M�馯���T$�B��J�3������@O�����M������T$�B��J�3������O�����M�����T$�B��J�3��`�����N�e����M�����T$�B�J�3��=�����N�B����M��j���T$�B�J�3�������N�����M��G���E����   �e���M�/��ËT$�B�J�3��������N������EЃ��   �e���M����ÍM������M������T$�BȋJ�3������hN�����M������M�����M�����M�����M���P���M�����T$�B��J�3��O����DN�T����M��|���T$�B��J�3��,���� N�1����M��Y���M��Q���M��I���M��aP���T$�B��J�3��������M������M��>P���M��6P���T$�B��J�3��������M������M��P���T$�B�J�3�������M�����M������M������M������T$�BȋJ�3��p�����M�u����M�����T$�B��J�3��M����lM�R����̋M��������M��}����T$�B�J�3�������R�"����̋E����   �e���M�8��ËT$�B��J�3��������K����������������̍M����T$�B��J�3������S����������������̍M���N���E܃��   �e���M��N��ËT$�B�J�3��o�����R�t������̍M���+���Eԃ��   �e���M��+��ËT$�B��J�3��/�����R�4������̍M��X���E����   �e���M�@��ËT$�B�J�3�������PR��������̍M��8N���E܃�t�e���M�$N��ËT$�B�J�3������tY�����M�� N���E܃�t�e���M��M��ËT$�B�J�3��{����PY�����M������M��pU���T$�BԋJ�3��P����,Y�U����M������M��EU���T$�B؋J�3��%����Y�*����M��b����M��U���Ẽ��   �e���M�r*��ËT$�BЋJ�3��������X������M������M���T���Ẽ��   �e���M�.*��ËT$�BЋJ�3�������X�����M�������M��T���T$�B؋J�3��r�����X�w����M������M��gT���T$�B؋J�3��G����xX�L����M������M��<T���T$�B̋J�3������TX�!����M��Y����M�T���T$�B��J�3�������0X������M��.����M���S���T$�BԋJ�3�������X������M������M��S���T$�B؋J�3�������W�����M�������M��S���T$�BԋJ�3��p�����W�u����M������M��eS���T$�B؋J�3��E�����W�J����M������M��:S���T$�BԋJ�3������|W�����M��W����M��S���T$�B؋J�3�������XW������M��,����M���R���T$�BԋJ�3�������4W������M������M��R���T$�B؋J�3������W�����M�������M��R���T$�BԋJ�3��n�����V�s����M������M��cR���T$�B؋J�3��C�����V�H����M������M��8R���T$�BԋJ�3�������V�����M��U����M��R���T$�B؋J�3��������V������M��*����M���Q���T$�BԋJ�3�������\V������M�������M��Q���T$�B؋J�3������8V�����M�������M��Q���T$�BԋJ�3��l����V�q����M������M��aQ���T$�B؋J�3��A�����U�F����M��~����M��6Q���T$�BԋJ�3�������U�����M��S����M��Q���T$�B؋J�3��������U������M��8I���M������T$�BċJ�3��������U������M��}����M������T$�B܋J�3������`U�����M��R����M�����T$�B܋J�3��j����<U�o�����������������̋E���t�e���M�|���ËT$�B��J�3��+����X]�0����M��X����M��P����T$�B��J�3�� ����4]�����M��-����E����   �e���M����ËT$�B�J�3�������]������M�������E����   �e���M�����ËT$�B�J�3�������\�����E���t�e���M��$��ËT$�B��J�3��X�����\�]����E���t�e���M�G��ËT$�B��J�3��(�����\�-����M��U����E����   �e���M�=���ËT$�B�J�3��������\������M������E����   �e���M����ËT$�B�J�3������\\�����M��$���Eԃ�t�e���M�����ËT$�B��J�3��x����8\�}����M������E����   �e���M����ËT$�B�J�3��<����\�A����M��F���M��q����Ẽ��   �e���M�iF��ËT$�BԋJ�3��������[������M��%����E����   �e���M����ËT$�B�J�3�������[������M�������E����   �e���M����ËT$�B�J�3�������[�����M���E���T$�B܋J�3��]�����[�b����Ẽ��   �e���M�z���ÍM��E���M��y����T$�BЋJ�3������`[�����Ẽ��   �e���M�6���ÍM��ME���M��5����T$�BЋJ�3�������<[������M��"E���M��
����T$�B؋J�3������[�����M���D���M��߾���T$�B؋J�3�������Z�����M���D���E܃�t�e���M�D��ËT$�B�J�3��G�����Z�L��������������̍M��D���T$�B�J�3�������]����������������̍M�8�����T����}4����L������   ��L�����M��O!��Ë�L������   ��L������X��������Ë�L������   ��L������h����!��Ë�L������   ��L�����M��� ��Ë�L������   ��L����M��� ��Ë�L����� �   ��L���ߍM�� ��ËT$��L�����H���3�������]���������������̍M��x ���T$�B��J�3��������_�����h�6j;h�r�E�P�����ËT$�B��J�3������\_�����M�������M�������EЃ��   �e���M�����ËT$�BЋJ�3��p����8_�u����M������M������EЃ��   �e���M�}���ÍM��t����T$�BЋJ�3��$����_�)����M��Q����M��I����EЃ��   �e���M�1���ÍM��(����M�� ����T$�BЋJ�3��������^������M�������M�������EЃ��   �e���M�����ÍM�������M�������M�������T$�BЋJ�3��t�����^�y����M������E����   �e���M�����ËE����   �e���M��p���ËT$�B��J�3�������^�$����M��L����E����   �e���M��4���ËE����   �e���M�����ËT$�B��J�3��������^�������������������̍M��H���E���   �e���M�H��ËT$�B��J�3�������`�����M��|H���E���   �e���M�dH��ËT$�B��J�3��C�����`�H����M��@H���E܃��   �e���M�(H��ËT$�B�J�3������``�����E����   �e���M�$���ÍM������T$�B�J�3�������<`������M�������E����   �e���M�����ËT$�B�J�3�������a�����M��̹���T$�B�J�3��l�����a�q����M�驹���E����   �e���M鑹��ËT$�B�J�3��0�����a�5����M����:m���T$�B��J�3��
�����a����h,7h�   h�r�E�P�����ËT$�B��J�3�������da������M����l���T$�B��J�3������@a�����M���>���M�������T$�BЋJ�3������a����������̍M�����T$�B��J�3��X���� b�]���������������̋M���������M��������T$�B��J�3������Tb������������������̋E܃��   �e���M�8���ÍM���E���T$�B��J�3��������b���������h!����Y����̃=�r uK�|r��t��rQ�@<�@�Ѓ��|r    V�5�r��t������V�j������r    ^�                                                                                                                                                           �f �f rf Vf Bf 2f "f �f     �d �d �d �d e e (e 4e Be Pe �d be pe ~e �e �e �e �e �e f |d rd fd ^d Td Jd Bd Xe ,d          !         ���            l; 0 �J�J�J�J�J�JKsrc/Commands.cpp    cmd-loadcontainer.tif   �; � �J�J� �J�J�JKcmd-preparecontainer.tif    Ocontainer.png  Ocontainer      GD&oMfP1MS),3SI %-3-ltru(zl(Th5w6/A::K,jI-7vNBU vO$FqmN-guAHc%ny)1r&wnyx62U 6qOMyfjBI9go$;Kblw93NwFX-kv9xq_GbHqkBKKCcY)0;R5BcYw:        �<` �"  !  1 �1 �$ �  �g �g �g �g 0! �g �g  h h  h ����@�0���Т�� �� �0�@�P�`�src/ContainerObject.cpp     333333�?ffffff�?      �?     �o@�<�9 ../../resource/_api/c4d_file.cpp    ../../resource/_api/c4d_file.cpp    res Progress Thread 0%  ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp %   ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ../../resource/_api/c4d_gui.cpp ~   |=�� �k �k �k  l l `l �l �l �l �l h=�� �{ �{  | |  | 0| @| P| �=�� �{ �{  | |  | 0| @| � �<�� �{ �{  | |  | 0| @| � >�� �{ �{  | |  | 0| @| @� �� �� �� о � �  � � 0� @� P� �� -DT�!	@      Y@     �f@     @�@�������������   %s  p:\applications\maxon\cinema 4d r13.061\resource\_api\c4d_general.h ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  ../../resource/_api/c4d_baseobject.cpp  `>0JpF�>pJ����MbP?res ../../resource/_api/c4d_resource.cpp    ../../resource/_api/c4d_resource.cpp    #   #   #   #   #   #   #   #   #   #   M_EDITOR    M_EDITOR    ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp  ../../resource/_api/c4d_basebitmap.cpp              �������?-DT�!�?      �-DT�!��               �       �../../resource/_api/c4d_pmain.cpp   ../../resource/_api/c4d_pmain.cpp   ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp    ../../resource/_api/c4d_basetime.cpp          �?   ����A  4&�kC �Ngm��C  4&�k�        ��������������(?`�������../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_libs/lib_ngon.cpp   ../../resource/_api/c4d_gv/ge_mtools.cpp    p?��?�� @��H@`��@��    �rsH                                                           `r�@�              ;;8;     p       ����    @    ;p        ����    @   T;           d;8;                4p�;           �;�;;8;    4p       ����    @   �;            Xp�;           �;�;;8;    Xp       ����    @   �;           <(<8;    �p       ����    @   <           T<d<(<8;    �p       ����    @   D<            �p�<           �<�<d<(<8;    �p       ����    @   �<            pT;            �p�<           ==4=    �p       ����    @   �<�p        ����    @   P=           `=4=                �pP=            q�=           �=�=    q        ����    @   �=            $q�=           �=�=4=    $q       ����    @   �=            @q$>           4>D>=4=    @q       ����    @   $>            \qt>           �>�>    \q        ����    @   t>           �>�>    tq        ����    @   �>            �q�>            ??�>    �q       ����    @   �>            �q<?           L?T?    �q        ����    @   <?            �q�?           �?�?    �q        ����    @   �?            �q�?           �?�?    �q        ����    @   �?            r@           $@,@    r        ����    @   @            $r\@           l@x@�>    $r       ����    @   \@            Hr�@           �@�@    Hr        ����    @   �@    �   i � � , X � �  X �  M x � � �  @ � �  X { � �  Y � �  X � *	 f	 �	 �	 
 W
 �
 �
 �
  & I t � � � ( K n � � � 
 - P s � �  a � � �  @ c � � � A � � � 5 ` � �  > i � � �  @ k � � �  B m � � �  D o � � �  F � � � ( X � �   8 t � � 0 S � �  1 i � � � � @ � � < � � 1 m � � ! D � � �   .  X  �  �                  ����@����Y   a"�   HC                       ����        "�   �C                       ����������   �"�   �C                       ���������       $"�   D                       "�   �C                       �����    �"�   dD                       "�   �D                       ����0    @   H   P    8���� ����"�   �D                       "�   <E                       �����    �   �   �   �   �   �    �   �   �	   �	   ����� "�   �E                       �����    �    �"�   �E                       ����P"�   F                       ����8    0"�   0F                       ��������������s������������������������p����M	    E	��������������|    t����?    7����'    �����    �    ����		    �   	    "	����7    '   /    P�����    �   �    ����8    (   0    Q�����    �   �    �����    �   �    �����k    [   c    �"�   �F                       "�   G                       "�   K                       "�   ,G                       "�   LG                       "�   �F                       "�   �F                       "�   lG                       "�   �G                       "�   dF                       "�   lF                       "�   tF                       "�   �F                       "�   �F                       "�   �G                       "�   �G                       "�   �F                       "�   |F                       "�   �F                       "�   �F                       "�   �F                       "�   �F                       �����    s   �   �   �   �    �"�   `K                       �����	    �	   �	   �	   �	   �	�����"�   �K                       ����[��������|���������k����H����%�������������f����C��������������A��������
�����	���������������    ������    ������    �����d    l�����
    �
�����
    �
�����
    �
����r
    z
����6
    O
����(    0   8�����        �����    �   ������    �   ����������             "�   �K                       "�   �L                       "�   �K                       "�   DL                       "�   ,M                       "�   �K                       "�   R                       "�   �L                       "�   TL                       "�   �K                       "�   �K                       "�   �K                       "�   �K                       "�   �K                       "�   dL                       "�   tL                       "�   �K                       "�   L                       "�   L                       "�   LM                       "�   L                       "�   L                       "�   M                       "�   �L                       "�   $L                       "�   ,L                       "�   �L                       "�   �L                       "�   �L                       "�   �L                       "�   �L                       "�   4L                       "�   <L                       ����1����9����A����I����Q   Y�����    �"�   @R                       ����h    `"�   tR                       ����(     "�   �R                       �����    �"�   �R                       �����"�   S                       ����6    >����    �����    ������    ������    �����_    g����4    <����	    �����    ������    ������    �����]    e����2    :����    �����    ������    ������    �����[    c����0    8����    �����    ������    ������    �����Y    a����.    6����{    �����P    X����     �����    ������    �   ������    �   �"�   <S                       "�   LS                       "�   \S                       "�   lS                       "�   |S                       "�   �S                       "�   �S                       "�   �S                       "�   �S                       "�   �S                       "�   �S                       "�   �S                       "�   �S                       "�   T                       "�   T                       "�   ,T                       "�   <T                       "�   LT                       "�   \T                       "�   lT                       "�   |T                       "�   �T                       "�   �T                       "�   �T                       "�   �T                       "�   U                       "�   $U                       "�   �T                       "�   �T                       "�   �T                       "�   �T                       ����K����s����C����p����T    L����!    )�����    �����    �����    �����[    S����#    �����    ������    �����    �����    ������    �   �����n    �   ������    �����������    �   �    �"�   �Y                       "�   �Y                       "�   �Y                       "�   hZ                       "�   �Z                       "�   �Y                       "�   �Y                       "�   �Y                       "�   �Z                       "�   Z                       "�   Z                       "�   (Z                       "�   8Z                       "�   �Y                       "�   �Y                       "�   HZ                       "�   XZ                       "�   �Z                       "�   �Y                       �����"�   |]                       "�   �]                       �����    �   �   �      6   U   t��������������������   �����W����_   x����'       ����k    [   c   �"�   ^                       "�   4^                       "�   �_                       "�   �_                       "�   d^                       "�   L^                       "�   ^                       "�   ^                       �����    �   �   �   �����    �      $   ,   4�����    ������    �����T    L����    "�   �_                       "�   `                       "�   `                       "�   ,`                       �������������������<���� ����& ����g    _����     "�   �`                       "�   �`                       "�   �`                       "�   �`                       "�   �`                       "�   �`                       "�   a                       ����P "�   b                       �����     � "�   Db                       �����     � "�   xb                           ����    ����    ����    ��    t�������    ����    ����    ��    ����    ����    ����    g�    ����    ����    ��������    ����    ����    ���������c         �d $0 �c         �f  0                     �f �f rf Vf Bf 2f "f �f     �d �d �d �d e e (e 4e Be Pe �d be pe ~e �e �e �e �e �e f |d rd fd ^d Td Jd Bd Xe ,d     x__CxxFrameHandler3  �free  malloc  ,memset  �floor 1_purecall (memcpy  k_libm_sse2_asin_precise m_libm_sse2_cos_precise  s_libm_sse2_sqrt_precise Q_CIfmod MSVCR110.dll  p ??1type_info@@UAE@XZ  s__CppXcptFilter _amsg_exit  �_malloc_crt �_initterm �_initterm_e 
_vsnprintf  |_lock �_unlock +_calloc_crt �__dllonexit "_onexit K_crt_debugger_hook  �__crtUnhandledException �__crtTerminateProcess ;?terminate@@YAXXZ �__clean_type_info_names_internal  p_except_handler4_common <EncodePointer DecodePointer �IsDebuggerPresent �IsProcessorFeaturePresent <QueryPerformanceCounter $GetCurrentProcessId (GetCurrentThreadId  �GetSystemTimeAsFileTime KERNEL32.dll      �n
R    g          g g g �� &g   containerobject.cdl c4d_main                                                                                                                                                                                                                  �:    .?AVCommandData@@   �:    .?AVBaseData@@  �:    .?AVLoadContainerCommand@@  �:    .?AVPrepareContainerCommand@@   x1�:    .?AVNodeData@@  �:    .?AVObjectData@@    �:    .?AVContainerObject@@   �:    .?AVSubDialog@@ �:    .?AVGeDialog@@  �:    .?AVGeUserArea@@    �:    .?AVGeModalDialog@@ �:    .?AViCustomGui@@    �:    .?AVNeighbor@@  �:    .?AVGeSortAndSearch@@   �:    .?AVDisjointNgonMesh@@  �:    .?AVC4DThread@@ �:    .?AVGeToolNode2D@@  �:    .?AVGeToolList2D@@  �:    .?AVGeToolDynArray@@    �:    .?AVGeToolDynArraySort@@    �:    .?AVtype_info@@ N�@���D        ����                                                                                                                                                                                                                                                                                                                                                                                                               �   0T0w0�0�01B1U1t1�142O2j2y2�2�2333F3�3�3�3g4�4�4�4�45"5@5�5�5�5�5%67)7<7N7]7z7�7�78$868=8f8o8�8�8�839D9V9`9�9�9�9�9":�:�:;e;�;�; <<0<a<�<�<�< ==@=l=�=�=�=�=�=>>/>Y>�>�>?c?q?�?�?�?      �   0060<0�031E1�12&2E2�2�2�2�23 3.3<3t3�3�3�3�34424G4a4q4C5V5j5�56*6]6}6�6�6*7D8H8L8P8T8X8\8`8d8s8�8�8�8$9R9z9�9�9:_:�:�:�:;A;�;<4<O<b<�<�<o=�=�=�=#>e>�>�>?g?�? 0    00&0b0~0�0�0�0R2�2�2�2�2�2
3 3%3B3~3�3�3�34"4^4�4�4�4�4�45A5q5�5�5�5�56M6u6�6�6�677l7�7�7 8(8A8a8�8�8�8�8�8�8�8Q9a9q9�9�9�9�9�9�9�9�9:!:5:S:a:y:�:�:�:�:�:;C;Q;i;w;�;�;�;�;�;<C<Q<i<<�<�<�<==.=D=^=n=�=�=�=�=>.>A>X>s>�>�>�>�>?!?8?S?�?�?�?�? @    10A0Q0q0�0�0�0�01!111S1a1{1�1�1�12!2A2a2q2�2�2�2�2�2�233!313A3Q3a3q3�3�3�3�3�3�3�3�3(4G4�4�4�4�45-5K5p5�5�516K6b6�6�6�6�67+7B7Y7p7�7�7�78)8@8�8�8�8�8�8�8�8919S9c9�9�9�9
::*:^:r:�:�:;1;V;v;�;�;�;<><`<~<�<�<=*=N=r=�=�=>>1>A>Q>a>�>�>�>�>�>�>�>??$?>?S?m?�?�?�?�?   P  d  010A0S0d0~0�0�0�0�0�031D1b1w1�1�1�1�12!212A2Q2a2q2�2�2�2�2�2�2313Q3a3q3�3�3�3�3�3�3�3�34!414N4q4�4�4�4�4�4�4�4�455!515A5Q5a5q5�5�5�5�5�5�5�566)6Q6q6�6�6�6�6�6�6�6�677!717A7q7�7�7�7�7�7�7�7�788#838U8v8�8�8�8�819A9Q9a9q9�9�9�9�9�9�9 ::2:c:t:�:�:�:�:�:;c;u;�;�;�;�;
< <A<[<�<�<�<�<=*=D=W=n=�=�=�=�=�=>">>>X>h>�>�>�>�>?!?1?a?�?�?�?�?�? `  �   0#0A0^0�0�0�0�0111A1Q1a1q1�1�1�1�1212`2�2�2�23+3a3�3�3�3�3�3�344!414A4Q4a4q4�4�4�4�4�4�4�4�455,5Q5a5�5�5�5�566A6d6z6�6�6�6�6�6V8]8d8k8r8y8�8�8�8�8�8�8�8�8�8�8�8S9g9�9�9�9�:r;�;�;<-<�<0=`=y=�=�=k>�>�>�>�>K?�?�?�?�? p  �   010Q0u0�0�0�01!1A1`1t1�1�1�1�1252U2q2�2�2�2�2 33(3F3j3�3�3�3�3�344=4e4�4�4�455a5�5�5�5!6A6a6�6�6�6757e7�7�7�78888�8�8�8�8%9Q9u9�9�9:#:=:N:�:5;a;�;�;�;�;�;Q<�<�<�=�=�=>3>C>�>�>�>!?A?a?�?�?�? �  �   %0U0q0�0�0C1T1v1�1�1�1�1232J2x2�2�2�23I3b3�3�3�34#4F4u4�4J5R5Z5v5�5Y6k6�6 7;7�78*828P8h88�8�8#939U9w9�9�9�9>:s:�:�:;h;�;�;<B<�<�<�<=O=�=�=�=>>'>i>�>�>!?z? �  �   0�0�0�0�01z1�12(2�2�2�233S3c3�304G4u4�445X5�5�5�5 6N6_6�6�6757s7�7�7�7�7#838i8�89#9�:�:�:�:X;3<C<}<�<�<�<=2=�=�=>M>}>�>�>?A?�?�?�? �  �   0_0�01_1�1�1O2�2�2?3�3�3/44�45_5�5�5A6�6�6(7�7�78a8�8�89M9�9�9�9+:M:}:�:�:;;>;�;�;><`<z<�<�<�<%=U=�=�=�=)>[>�>�>?=?a?�?�?�? �  �   !0Q0�0�0�0!1C1S1t1�12-2d2�2�2�2_3�3�3�3�34$4v4�4�4�4�45555k5�5�5�56-6X6n6�6�6�6�677B7e7�7�7'8�89�9�9�9�9�9�9 ::::.:!;�;�;�;�;�;�;�;�;�;v<{<�<�<�<�<�<)=s=�=�=�=�=�=�=	>A>o>�?�?   �  �   0C0R0�01#1X1�1�1�1!2E2q2�2�2�2�2�2�23C3V3p3�3�3�3�3
44.4G4u4�4�4�4�4!515A5�5�5�5�5�56:6Z6t6�6�6797Y7}7�7�78+8C8�8�8�8�899Q9�9�9�9�9�9�9P:g:~:�:�:;);[;`;x;�;�;�;+<Y<�<�<=s=�=�=>>4>9>N>{>�>�>�>�>?"?~?�?�? �  �   /0N0|0�0�0�0�061N1e1|1�1�1�1�1292\2�2�2�2!3�3�34�4�4�4456.6�67�7�78c8s8�8�89�9�9�9:*:J:�:�:�:�:S<`<�<�<�<==0=�=�=�=>$>B>^>x>�>�>�>??G?a?�?�?�?�?�?   �  �   0000�0�0�0�0151Q1u1�1�1�12!2A2a2q2�2�2�2�2�2�2�2�23!313Q3q3�3�3�3�34 4�4�4545s5�5�536D6�6�6C7T7�78S8c8w8�839C9W9�9:$:�:�:;#;�;�;�;i<�<�<�<K=�=�=>1>O>m>�>�>�>W?�?�?   �  �   &0A0_0}0�0�0�0g1�1�1#242�2�2�23S3c3w3�334D4�4�4�45c5s5�56C6T6�6�637C7�7�78�8�8�8�8#939G9�9::�:�:�:;{;�;�;I<d<�<�<+=�=�=�=�=>!>E>c>u>�>�>?4?R?�?�?�?�?�?   (  0a0�0�0�0�01!111Q1q1�1�1�1%2Q2a2q2�2�2�2�2�2�2�2 33
33'3Q3a3q3�3�3�3�3�3414a4q4�4�4�45>5z5�5�5-6^6�6�677!7�7�7�7�7858a8q8�8�8�8�89A9e9�9�9�9�9:A:Q:a:q:�:�:�:�:;;!;1;A;Q;a;q;�;�;�;�;�;�;	<,<C<U<�<�<�<�<�<�<= =c=t=�=�=�=�=>!>1>A>Q>a>q>�>�>�>�>�>�>�>�>??!?1?C?Q??�?�?�?�?      00!0O0�0�0�011Q1a1q1�1�1�1�1�1�1�1�122#242R2j2�2�2�2�23343D3�3�3�3�3414A4Q4a4q4�4�4�4�4�4�4A5Q5a5q5�5�5�5�5�5�5D6�6�6�6757a7�7�7�7�78!8T8o8�8�89=9`9�9�9�9�9�9:(:B:R:�:�:�:�:;S;b;t;�;�;�;3<D<^<r<�<�<�<==s=�=�=�=�=#>9>N>^>�>�>�>?B?X?�?�?�?�?     20H0�0�0�0�0�011!111A1Q1a1q1�1�1�1�1�1�1�1 2a2q2�2�2�2�2�2�2�2�233!313A3Q3a3q3�3�3�34!4A4a4�4�4�4�45!5X5�5�5�56!6E6s6�6�6�6�67<7�7�7�78!818e8~8�8�8�8929X9k9�9�9�9	:,:=:e:�:�:�:�:;1;Q;q;�;�;<!<Q<�<�<�<=1=Q=q=�=�=�=�=>A>x>�>�>�>�>?1?Q?q?�?�?�? 0 �   0=0Q0f0�0P1�1�12,2R2�2�2�2�23D3�3�3�34!4A4a4�4�4�4�45!5E5q5�5�5�5�5616U6�6�6�6�677$7A7q7�7�78a8�8�8�8�89K9�9�9�9:D:b:�:�:�:�:;*;K;<!<f<n<�<�<�<4=E? @ �   262~2�2�2�23_3x35 5$5(5;5a5q5�5�5�5�5B6U6Z6q6�6�6�6A7Q7d7�7�7`8�8�8�8�859�9�9�9�98:=:�:�;�;�;�;�;�;�;�;�;C<X<�<�<�<=c>?�?�? P    0c0q0�0�0�0;1c1�1�122C2T2o2y2�2�2�2�2�2�2�2383R3�3�3�3�34$4?4I4U4h44�4�4�4�4�45"5g5�5�5�5�5�5�56<6N6b6�6�6�6�6�6�67"7<7O7Z7~7�7�7�78&898D8h8�8�8�8�8�8�8 9:9\9y9�9�9�9�9::%:8:O:b:|:�:�:�:�:�:7;T;f;y;�;�;�;�;<<1<<<`<z<�<�<�<�<�<='=I=f=x=�=�=�=T>i>�>�>�>�>?"?*?A?�?�? ` �   0N0w0�0�011*121I1�1�12P2y2�2�23"3+343F3Q3k324b4�4�4�4B5f5�5�5�5"6J6s6�6�6727b7�7�7�78R8�8�8�89L9r9�9�9�9A:i:�:�:�:�:�:;@;h;�;�;<<%<x<�<�<A={=�=>B>�>�>�>"?b?�?�? p �   "0R0�0�01R1�1�1�1"2b2�2�23#373�3�34b4�4�425r5�56B6�6�677&7I7�7�7�7�78!818a8�8�8�89%9Q9q9�9�9�9�9�9:A:a:�:�:�:�:�:�:;;E;u;�;�;�;<#<3<E<b<{<�<�<�<=%=U=�=�=�=�=>A>a>�>�>�>�>?!?A?c?s?�?�?�? � d   !010U0�0�0�0�0q1�1�1�112A2Q2q2�2�2C3Q3)4S4`4r4|4�4�4A5�5�56E7q7�7�7�7�7�9�9
::7:b:=;V;�<> � 4   �6�7�7&9�9�;�;�;�;�;�;�;0<E<�<�<d=�=F>=?U?   � �   �02q3�34&4<4e4�4�4�4�4�4�4�4�5�8:9B9K9W9q9�9:a:�:�:�:A;q;�;�;�;�;<<5<n<�<�<�<�<�<�<�<�<�<�<�<==I=�=�=+>s>�>�>�>�>�>?$?c?q?�?�?�?�?�? � �   
00"070_0p0u0�01.1Q1n1�1�1�1D2J2V2_2f2�2�2�2�2�2*383m3�3�3�3�3�3�3Q4k4�4�4�4�45!515A5i5p5�5�5�5616Q6q6�6�6�6�67!7A7a7�7�7�7�78!8A8a8�8�8�8�89!9A9a9�9�9�9!:a:�:�:�:;!;A;a;�;�;�;�;<!<D<�<�<�<=!=A=a=�=�=�=�=>!>E>a>�>�>�>�>?!?U?�?�? � @   30�0�0�7�7�7�73888U8Z8>9C9w9|9F:K:{:�:>;C;y;~;�;�;%>P>   � <   �3�3 4444|6�6�6:�<�<=B=�=�=>B>�>�>�>"?b?�?�?�? � \   20b0�0�0�0"1R1�1�12R2�2�23R3�3�324�4�45B5�5W78	8#8c8q8�8�8�8�:;	; <P<�>�>g?l?�? � @  0�0�0�0�0151e1�1�1�12w2�2�2�3�3�3
4!454e4�4�4�4�455u5�5�5616Q6e6�6�6�6�6(72777<7R7^77�7�7�7�7�7�7�788%8/858=8m8u8z88�8�8�8�8�8�8�8999.969M9S9�9�9�9�9-:_:�:�:�:�:�:�:�:�:�:�:;; ;3;H;S;i;�;�;�;�;�;�;�;�;�;5<;<A<G<M<S<Z<a<h<o<v<}<�<�<�<�<�<�<�<�<�<�<�<�< =	==�=�=�=�=V>[>m>�>�>�>H?k?w?�?�?�?�?�?�?�?     �    00 0&0+0A0^0�0�0�0�0�0�0�0�0�0�0�0�0*1A1H1{1�1�1�12>2j2�2�2�2�23j3�3"4_4�4�4�4�45R5�5�5.6j6�6�6�67k7�7�78j8�8<9x9�9
:-:i:�:�:�:;8;[;�;�;�;�;:<]<�<�<�<�<=?=b=�=�=�=(>s>�>�>�>?R?u?�?�?  �   
0S0�0�01G1r1�1�1%2P2{2�2�2�2'3R3}3�3�3�3)4T44�4�4 5+5V5�5�5�56-6X6�6�6�6:7j7�7�78J8�8�89B9e9�9�9:C:{:�:�;�;�;�;<R<�<�<N=�=�=C>>�>�>3?V?�?�?�?�?�?         0@0j0�0�0111$161A1[1 0   �0�0�0�0�0�0�0�0�0�0�0�0�0111 1$1(1,1014181 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�24444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555T6X6\6`6d69999 9�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;4;8;P;`;d;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;<<< <(<@<P<T<X<\<d<|<�<�<�<�<�<�<�<�<�<�<�<�<�<====0=4=L=\=`=t=x=�=�=�=�=�=�=�=�=�=�=�=�=>> >0>4>8><>D>\>l>p>�>�>�>�>�>�>�>�>�>�>�> ???$?4?8?H?L?T?l?|?�?�?�?�?�?�?�?�?�?�?�? @ �  00 0$0,0D0T0X0h0l0p0x0�0�0�0�0�0�0�0L3T3\3h3�3�3�3�3�3�3�3�3 4444$4H4h4p4|4�4�4�4�4�4�4�4�4�4 5@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�56646<6H6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78<8`8�8�8�8�8989\9�9�9�9�9:4:X:|:�:�:�:;;; ;(;0;8;D;d;l;t;|;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ==== =(=0=8=@=H=P=X=`=h=t=�=�=�=>(>L>p>�>�>�> ?$?H?l?�?�?�?�?   P �   0D0h0�0�0�0�01@1d1�1�1�1�122$2,242<2D2L2X2x2�2�2�2�2�2�2�2�23 3@3H3P3X3`3h3p3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585D5h5�5�5�5�56@6d6�6�6�6�67<7`7�7�7�7�7888\8�8�8�8�8949X9|9�9�9�9�9�9�9�9�9�9�9�9�9�9::::$:,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�: ;D;h;�;�;�;�;<@<d<�<�<�<�<=<=`=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>H>P>X>`>h>p>x>�>�>�>�>�>?@?d?�?�?�?�?�?�?�?�?�?�?�?�? ` d    0000 0(00080D0h0�0�0�0�0�0�0�0�0 1111$1H1l1�1�1�1�12(2H2P2\2|2�2�2�2�2�2�23,303L3P3 p 4    0040X0�0�0�0�0�0�01$1@1\1t1�1�1�1�12$2H2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                